magic
tech sky130A
magscale 1 2
timestamp 1659965804
<< nwell >>
rect 1066 129733 129758 130299
rect 1066 128645 129758 129211
rect 1066 127557 129758 128123
rect 1066 126469 129758 127035
rect 1066 125381 129758 125947
rect 1066 124293 129758 124859
rect 1066 123205 129758 123771
rect 1066 122117 129758 122683
rect 1066 121029 129758 121595
rect 1066 119941 129758 120507
rect 1066 118853 129758 119419
rect 1066 117765 129758 118331
rect 1066 116677 129758 117243
rect 1066 115589 129758 116155
rect 1066 114501 129758 115067
rect 1066 113413 129758 113979
rect 1066 112325 129758 112891
rect 1066 111237 129758 111803
rect 1066 110149 129758 110715
rect 1066 109061 129758 109627
rect 1066 107973 129758 108539
rect 1066 106885 129758 107451
rect 1066 105797 129758 106363
rect 1066 104709 129758 105275
rect 1066 103621 129758 104187
rect 1066 102533 129758 103099
rect 1066 101445 129758 102011
rect 1066 100357 129758 100923
rect 1066 99269 129758 99835
rect 1066 98181 129758 98747
rect 1066 97093 129758 97659
rect 1066 96005 129758 96571
rect 1066 94917 129758 95483
rect 1066 93829 129758 94395
rect 1066 92741 129758 93307
rect 1066 91653 129758 92219
rect 1066 90565 129758 91131
rect 1066 89477 129758 90043
rect 1066 88389 129758 88955
rect 1066 87301 129758 87867
rect 1066 86213 129758 86779
rect 1066 85125 129758 85691
rect 1066 84037 129758 84603
rect 1066 82949 129758 83515
rect 1066 81861 129758 82427
rect 1066 80773 129758 81339
rect 1066 79685 129758 80251
rect 1066 78597 129758 79163
rect 1066 77509 129758 78075
rect 1066 76421 129758 76987
rect 1066 75333 129758 75899
rect 1066 74245 129758 74811
rect 1066 73157 129758 73723
rect 1066 72069 129758 72635
rect 1066 70981 129758 71547
rect 1066 69893 129758 70459
rect 1066 68805 129758 69371
rect 1066 67717 129758 68283
rect 1066 66629 129758 67195
rect 1066 65541 129758 66107
rect 1066 64453 129758 65019
rect 1066 63365 129758 63931
rect 1066 62277 129758 62843
rect 1066 61189 129758 61755
rect 1066 60101 129758 60667
rect 1066 59013 129758 59579
rect 1066 57925 129758 58491
rect 1066 56837 129758 57403
rect 1066 55749 129758 56315
rect 1066 54661 129758 55227
rect 1066 53573 129758 54139
rect 1066 52485 129758 53051
rect 1066 51397 129758 51963
rect 1066 50309 129758 50875
rect 1066 49221 129758 49787
rect 1066 48133 129758 48699
rect 1066 47045 129758 47611
rect 1066 45957 129758 46523
rect 1066 44869 129758 45435
rect 1066 43781 129758 44347
rect 1066 42693 129758 43259
rect 1066 41605 129758 42171
rect 1066 40517 129758 41083
rect 1066 39429 129758 39995
rect 1066 38341 129758 38907
rect 1066 37253 129758 37819
rect 1066 36165 129758 36731
rect 1066 35077 129758 35643
rect 1066 33989 129758 34555
rect 1066 32901 129758 33467
rect 1066 31813 129758 32379
rect 1066 30725 129758 31291
rect 1066 29637 129758 30203
rect 1066 28549 129758 29115
rect 1066 27461 129758 28027
rect 1066 26373 129758 26939
rect 1066 25285 129758 25851
rect 1066 24197 129758 24763
rect 1066 23109 129758 23675
rect 1066 22021 129758 22587
rect 1066 20933 129758 21499
rect 1066 19845 129758 20411
rect 1066 18757 129758 19323
rect 1066 17669 129758 18235
rect 1066 16581 129758 17147
rect 1066 15493 129758 16059
rect 1066 14405 129758 14971
rect 1066 13317 129758 13883
rect 1066 12229 129758 12795
rect 1066 11141 129758 11707
rect 1066 10053 129758 10619
rect 1066 8965 129758 9531
rect 1066 7877 129758 8443
rect 1066 6789 129758 7355
rect 1066 5701 129758 6267
rect 1066 4613 129758 5179
rect 1066 3525 129758 4091
rect 1066 2437 129758 3003
<< obsli1 >>
rect 1104 2159 129720 130577
<< obsm1 >>
rect 1104 484 129720 131572
<< metal2 >>
rect 3606 132223 3662 133023
rect 4342 132223 4398 133023
rect 5078 132223 5134 133023
rect 5814 132223 5870 133023
rect 6550 132223 6606 133023
rect 7286 132223 7342 133023
rect 8022 132223 8078 133023
rect 8758 132223 8814 133023
rect 9494 132223 9550 133023
rect 10230 132223 10286 133023
rect 10966 132223 11022 133023
rect 11702 132223 11758 133023
rect 12438 132223 12494 133023
rect 13174 132223 13230 133023
rect 13910 132223 13966 133023
rect 14646 132223 14702 133023
rect 15382 132223 15438 133023
rect 16118 132223 16174 133023
rect 16854 132223 16910 133023
rect 17590 132223 17646 133023
rect 18326 132223 18382 133023
rect 19062 132223 19118 133023
rect 19798 132223 19854 133023
rect 20534 132223 20590 133023
rect 21270 132223 21326 133023
rect 22006 132223 22062 133023
rect 22742 132223 22798 133023
rect 23478 132223 23534 133023
rect 24214 132223 24270 133023
rect 24950 132223 25006 133023
rect 25686 132223 25742 133023
rect 26422 132223 26478 133023
rect 27158 132223 27214 133023
rect 27894 132223 27950 133023
rect 28630 132223 28686 133023
rect 29366 132223 29422 133023
rect 30102 132223 30158 133023
rect 30838 132223 30894 133023
rect 31574 132223 31630 133023
rect 32310 132223 32366 133023
rect 33046 132223 33102 133023
rect 33782 132223 33838 133023
rect 34518 132223 34574 133023
rect 35254 132223 35310 133023
rect 35990 132223 36046 133023
rect 36726 132223 36782 133023
rect 37462 132223 37518 133023
rect 38198 132223 38254 133023
rect 38934 132223 38990 133023
rect 39670 132223 39726 133023
rect 40406 132223 40462 133023
rect 41142 132223 41198 133023
rect 41878 132223 41934 133023
rect 42614 132223 42670 133023
rect 43350 132223 43406 133023
rect 44086 132223 44142 133023
rect 44822 132223 44878 133023
rect 45558 132223 45614 133023
rect 46294 132223 46350 133023
rect 47030 132223 47086 133023
rect 47766 132223 47822 133023
rect 48502 132223 48558 133023
rect 49238 132223 49294 133023
rect 49974 132223 50030 133023
rect 50710 132223 50766 133023
rect 51446 132223 51502 133023
rect 52182 132223 52238 133023
rect 52918 132223 52974 133023
rect 53654 132223 53710 133023
rect 54390 132223 54446 133023
rect 55126 132223 55182 133023
rect 55862 132223 55918 133023
rect 56598 132223 56654 133023
rect 57334 132223 57390 133023
rect 58070 132223 58126 133023
rect 58806 132223 58862 133023
rect 59542 132223 59598 133023
rect 60278 132223 60334 133023
rect 61014 132223 61070 133023
rect 61750 132223 61806 133023
rect 62486 132223 62542 133023
rect 63222 132223 63278 133023
rect 63958 132223 64014 133023
rect 64694 132223 64750 133023
rect 65430 132223 65486 133023
rect 66166 132223 66222 133023
rect 66902 132223 66958 133023
rect 67638 132223 67694 133023
rect 68374 132223 68430 133023
rect 69110 132223 69166 133023
rect 69846 132223 69902 133023
rect 70582 132223 70638 133023
rect 71318 132223 71374 133023
rect 72054 132223 72110 133023
rect 72790 132223 72846 133023
rect 73526 132223 73582 133023
rect 74262 132223 74318 133023
rect 74998 132223 75054 133023
rect 75734 132223 75790 133023
rect 76470 132223 76526 133023
rect 77206 132223 77262 133023
rect 77942 132223 77998 133023
rect 78678 132223 78734 133023
rect 79414 132223 79470 133023
rect 80150 132223 80206 133023
rect 80886 132223 80942 133023
rect 81622 132223 81678 133023
rect 82358 132223 82414 133023
rect 83094 132223 83150 133023
rect 83830 132223 83886 133023
rect 84566 132223 84622 133023
rect 85302 132223 85358 133023
rect 86038 132223 86094 133023
rect 86774 132223 86830 133023
rect 87510 132223 87566 133023
rect 88246 132223 88302 133023
rect 88982 132223 89038 133023
rect 89718 132223 89774 133023
rect 90454 132223 90510 133023
rect 91190 132223 91246 133023
rect 91926 132223 91982 133023
rect 92662 132223 92718 133023
rect 93398 132223 93454 133023
rect 94134 132223 94190 133023
rect 94870 132223 94926 133023
rect 95606 132223 95662 133023
rect 96342 132223 96398 133023
rect 97078 132223 97134 133023
rect 97814 132223 97870 133023
rect 98550 132223 98606 133023
rect 99286 132223 99342 133023
rect 100022 132223 100078 133023
rect 100758 132223 100814 133023
rect 101494 132223 101550 133023
rect 102230 132223 102286 133023
rect 102966 132223 103022 133023
rect 103702 132223 103758 133023
rect 104438 132223 104494 133023
rect 105174 132223 105230 133023
rect 105910 132223 105966 133023
rect 106646 132223 106702 133023
rect 107382 132223 107438 133023
rect 108118 132223 108174 133023
rect 108854 132223 108910 133023
rect 109590 132223 109646 133023
rect 110326 132223 110382 133023
rect 111062 132223 111118 133023
rect 111798 132223 111854 133023
rect 112534 132223 112590 133023
rect 113270 132223 113326 133023
rect 114006 132223 114062 133023
rect 114742 132223 114798 133023
rect 115478 132223 115534 133023
rect 116214 132223 116270 133023
rect 116950 132223 117006 133023
rect 117686 132223 117742 133023
rect 118422 132223 118478 133023
rect 119158 132223 119214 133023
rect 119894 132223 119950 133023
rect 120630 132223 120686 133023
rect 121366 132223 121422 133023
rect 122102 132223 122158 133023
rect 122838 132223 122894 133023
rect 123574 132223 123630 133023
rect 124310 132223 124366 133023
rect 125046 132223 125102 133023
rect 125782 132223 125838 133023
rect 126518 132223 126574 133023
rect 127254 132223 127310 133023
rect 10046 0 10102 800
rect 10230 0 10286 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 10966 0 11022 800
rect 11150 0 11206 800
rect 11334 0 11390 800
rect 11518 0 11574 800
rect 11702 0 11758 800
rect 11886 0 11942 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12806 0 12862 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13358 0 13414 800
rect 13542 0 13598 800
rect 13726 0 13782 800
rect 13910 0 13966 800
rect 14094 0 14150 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14646 0 14702 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15198 0 15254 800
rect 15382 0 15438 800
rect 15566 0 15622 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16670 0 16726 800
rect 16854 0 16910 800
rect 17038 0 17094 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18878 0 18934 800
rect 19062 0 19118 800
rect 19246 0 19302 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20534 0 20590 800
rect 20718 0 20774 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21270 0 21326 800
rect 21454 0 21510 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22374 0 22430 800
rect 22558 0 22614 800
rect 22742 0 22798 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23294 0 23350 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23846 0 23902 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24766 0 24822 800
rect 24950 0 25006 800
rect 25134 0 25190 800
rect 25318 0 25374 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26238 0 26294 800
rect 26422 0 26478 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 26974 0 27030 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28262 0 28318 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28814 0 28870 800
rect 28998 0 29054 800
rect 29182 0 29238 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30654 0 30710 800
rect 30838 0 30894 800
rect 31022 0 31078 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32126 0 32182 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32678 0 32734 800
rect 32862 0 32918 800
rect 33046 0 33102 800
rect 33230 0 33286 800
rect 33414 0 33470 800
rect 33598 0 33654 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34150 0 34206 800
rect 34334 0 34390 800
rect 34518 0 34574 800
rect 34702 0 34758 800
rect 34886 0 34942 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35438 0 35494 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 35990 0 36046 800
rect 36174 0 36230 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36726 0 36782 800
rect 36910 0 36966 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 38014 0 38070 800
rect 38198 0 38254 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39854 0 39910 800
rect 40038 0 40094 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40590 0 40646 800
rect 40774 0 40830 800
rect 40958 0 41014 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41878 0 41934 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42430 0 42486 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 42982 0 43038 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43718 0 43774 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44454 0 44510 800
rect 44638 0 44694 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45558 0 45614 800
rect 45742 0 45798 800
rect 45926 0 45982 800
rect 46110 0 46166 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46662 0 46718 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47582 0 47638 800
rect 47766 0 47822 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49606 0 49662 800
rect 49790 0 49846 800
rect 49974 0 50030 800
rect 50158 0 50214 800
rect 50342 0 50398 800
rect 50526 0 50582 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51630 0 51686 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52182 0 52238 800
rect 52366 0 52422 800
rect 52550 0 52606 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54574 0 54630 800
rect 54758 0 54814 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55310 0 55366 800
rect 55494 0 55550 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56230 0 56286 800
rect 56414 0 56470 800
rect 56598 0 56654 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57150 0 57206 800
rect 57334 0 57390 800
rect 57518 0 57574 800
rect 57702 0 57758 800
rect 57886 0 57942 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58438 0 58494 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59358 0 59414 800
rect 59542 0 59598 800
rect 59726 0 59782 800
rect 59910 0 59966 800
rect 60094 0 60150 800
rect 60278 0 60334 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60830 0 60886 800
rect 61014 0 61070 800
rect 61198 0 61254 800
rect 61382 0 61438 800
rect 61566 0 61622 800
rect 61750 0 61806 800
rect 61934 0 61990 800
rect 62118 0 62174 800
rect 62302 0 62358 800
rect 62486 0 62542 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63406 0 63462 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 63958 0 64014 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64694 0 64750 800
rect 64878 0 64934 800
rect 65062 0 65118 800
rect 65246 0 65302 800
rect 65430 0 65486 800
rect 65614 0 65670 800
rect 65798 0 65854 800
rect 65982 0 66038 800
rect 66166 0 66222 800
rect 66350 0 66406 800
rect 66534 0 66590 800
rect 66718 0 66774 800
rect 66902 0 66958 800
rect 67086 0 67142 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67638 0 67694 800
rect 67822 0 67878 800
rect 68006 0 68062 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68742 0 68798 800
rect 68926 0 68982 800
rect 69110 0 69166 800
rect 69294 0 69350 800
rect 69478 0 69534 800
rect 69662 0 69718 800
rect 69846 0 69902 800
rect 70030 0 70086 800
rect 70214 0 70270 800
rect 70398 0 70454 800
rect 70582 0 70638 800
rect 70766 0 70822 800
rect 70950 0 71006 800
rect 71134 0 71190 800
rect 71318 0 71374 800
rect 71502 0 71558 800
rect 71686 0 71742 800
rect 71870 0 71926 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72422 0 72478 800
rect 72606 0 72662 800
rect 72790 0 72846 800
rect 72974 0 73030 800
rect 73158 0 73214 800
rect 73342 0 73398 800
rect 73526 0 73582 800
rect 73710 0 73766 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74262 0 74318 800
rect 74446 0 74502 800
rect 74630 0 74686 800
rect 74814 0 74870 800
rect 74998 0 75054 800
rect 75182 0 75238 800
rect 75366 0 75422 800
rect 75550 0 75606 800
rect 75734 0 75790 800
rect 75918 0 75974 800
rect 76102 0 76158 800
rect 76286 0 76342 800
rect 76470 0 76526 800
rect 76654 0 76710 800
rect 76838 0 76894 800
rect 77022 0 77078 800
rect 77206 0 77262 800
rect 77390 0 77446 800
rect 77574 0 77630 800
rect 77758 0 77814 800
rect 77942 0 77998 800
rect 78126 0 78182 800
rect 78310 0 78366 800
rect 78494 0 78550 800
rect 78678 0 78734 800
rect 78862 0 78918 800
rect 79046 0 79102 800
rect 79230 0 79286 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80150 0 80206 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80702 0 80758 800
rect 80886 0 80942 800
rect 81070 0 81126 800
rect 81254 0 81310 800
rect 81438 0 81494 800
rect 81622 0 81678 800
rect 81806 0 81862 800
rect 81990 0 82046 800
rect 82174 0 82230 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82726 0 82782 800
rect 82910 0 82966 800
rect 83094 0 83150 800
rect 83278 0 83334 800
rect 83462 0 83518 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84014 0 84070 800
rect 84198 0 84254 800
rect 84382 0 84438 800
rect 84566 0 84622 800
rect 84750 0 84806 800
rect 84934 0 84990 800
rect 85118 0 85174 800
rect 85302 0 85358 800
rect 85486 0 85542 800
rect 85670 0 85726 800
rect 85854 0 85910 800
rect 86038 0 86094 800
rect 86222 0 86278 800
rect 86406 0 86462 800
rect 86590 0 86646 800
rect 86774 0 86830 800
rect 86958 0 87014 800
rect 87142 0 87198 800
rect 87326 0 87382 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88062 0 88118 800
rect 88246 0 88302 800
rect 88430 0 88486 800
rect 88614 0 88670 800
rect 88798 0 88854 800
rect 88982 0 89038 800
rect 89166 0 89222 800
rect 89350 0 89406 800
rect 89534 0 89590 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90086 0 90142 800
rect 90270 0 90326 800
rect 90454 0 90510 800
rect 90638 0 90694 800
rect 90822 0 90878 800
rect 91006 0 91062 800
rect 91190 0 91246 800
rect 91374 0 91430 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 91926 0 91982 800
rect 92110 0 92166 800
rect 92294 0 92350 800
rect 92478 0 92534 800
rect 92662 0 92718 800
rect 92846 0 92902 800
rect 93030 0 93086 800
rect 93214 0 93270 800
rect 93398 0 93454 800
rect 93582 0 93638 800
rect 93766 0 93822 800
rect 93950 0 94006 800
rect 94134 0 94190 800
rect 94318 0 94374 800
rect 94502 0 94558 800
rect 94686 0 94742 800
rect 94870 0 94926 800
rect 95054 0 95110 800
rect 95238 0 95294 800
rect 95422 0 95478 800
rect 95606 0 95662 800
rect 95790 0 95846 800
rect 95974 0 96030 800
rect 96158 0 96214 800
rect 96342 0 96398 800
rect 96526 0 96582 800
rect 96710 0 96766 800
rect 96894 0 96950 800
rect 97078 0 97134 800
rect 97262 0 97318 800
rect 97446 0 97502 800
rect 97630 0 97686 800
rect 97814 0 97870 800
rect 97998 0 98054 800
rect 98182 0 98238 800
rect 98366 0 98422 800
rect 98550 0 98606 800
rect 98734 0 98790 800
rect 98918 0 98974 800
rect 99102 0 99158 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99654 0 99710 800
rect 99838 0 99894 800
rect 100022 0 100078 800
rect 100206 0 100262 800
rect 100390 0 100446 800
rect 100574 0 100630 800
rect 100758 0 100814 800
rect 100942 0 100998 800
rect 101126 0 101182 800
rect 101310 0 101366 800
rect 101494 0 101550 800
rect 101678 0 101734 800
rect 101862 0 101918 800
rect 102046 0 102102 800
rect 102230 0 102286 800
rect 102414 0 102470 800
rect 102598 0 102654 800
rect 102782 0 102838 800
rect 102966 0 103022 800
rect 103150 0 103206 800
rect 103334 0 103390 800
rect 103518 0 103574 800
rect 103702 0 103758 800
rect 103886 0 103942 800
rect 104070 0 104126 800
rect 104254 0 104310 800
rect 104438 0 104494 800
rect 104622 0 104678 800
rect 104806 0 104862 800
rect 104990 0 105046 800
rect 105174 0 105230 800
rect 105358 0 105414 800
rect 105542 0 105598 800
rect 105726 0 105782 800
rect 105910 0 105966 800
rect 106094 0 106150 800
rect 106278 0 106334 800
rect 106462 0 106518 800
rect 106646 0 106702 800
rect 106830 0 106886 800
rect 107014 0 107070 800
rect 107198 0 107254 800
rect 107382 0 107438 800
rect 107566 0 107622 800
rect 107750 0 107806 800
rect 107934 0 107990 800
rect 108118 0 108174 800
rect 108302 0 108358 800
rect 108486 0 108542 800
rect 108670 0 108726 800
rect 108854 0 108910 800
rect 109038 0 109094 800
rect 109222 0 109278 800
rect 109406 0 109462 800
rect 109590 0 109646 800
rect 109774 0 109830 800
rect 109958 0 110014 800
rect 110142 0 110198 800
rect 110326 0 110382 800
rect 110510 0 110566 800
rect 110694 0 110750 800
rect 110878 0 110934 800
rect 111062 0 111118 800
rect 111246 0 111302 800
rect 111430 0 111486 800
rect 111614 0 111670 800
rect 111798 0 111854 800
rect 111982 0 112038 800
rect 112166 0 112222 800
rect 112350 0 112406 800
rect 112534 0 112590 800
rect 112718 0 112774 800
rect 112902 0 112958 800
rect 113086 0 113142 800
rect 113270 0 113326 800
rect 113454 0 113510 800
rect 113638 0 113694 800
rect 113822 0 113878 800
rect 114006 0 114062 800
rect 114190 0 114246 800
rect 114374 0 114430 800
rect 114558 0 114614 800
rect 114742 0 114798 800
rect 114926 0 114982 800
rect 115110 0 115166 800
rect 115294 0 115350 800
rect 115478 0 115534 800
rect 115662 0 115718 800
rect 115846 0 115902 800
rect 116030 0 116086 800
rect 116214 0 116270 800
rect 116398 0 116454 800
rect 116582 0 116638 800
rect 116766 0 116822 800
rect 116950 0 117006 800
rect 117134 0 117190 800
rect 117318 0 117374 800
rect 117502 0 117558 800
rect 117686 0 117742 800
rect 117870 0 117926 800
rect 118054 0 118110 800
rect 118238 0 118294 800
rect 118422 0 118478 800
rect 118606 0 118662 800
rect 118790 0 118846 800
rect 118974 0 119030 800
rect 119158 0 119214 800
rect 119342 0 119398 800
rect 119526 0 119582 800
rect 119710 0 119766 800
rect 119894 0 119950 800
rect 120078 0 120134 800
rect 120262 0 120318 800
rect 120446 0 120502 800
rect 120630 0 120686 800
rect 120814 0 120870 800
<< obsm2 >>
rect 1122 132167 3550 132274
rect 3718 132167 4286 132274
rect 4454 132167 5022 132274
rect 5190 132167 5758 132274
rect 5926 132167 6494 132274
rect 6662 132167 7230 132274
rect 7398 132167 7966 132274
rect 8134 132167 8702 132274
rect 8870 132167 9438 132274
rect 9606 132167 10174 132274
rect 10342 132167 10910 132274
rect 11078 132167 11646 132274
rect 11814 132167 12382 132274
rect 12550 132167 13118 132274
rect 13286 132167 13854 132274
rect 14022 132167 14590 132274
rect 14758 132167 15326 132274
rect 15494 132167 16062 132274
rect 16230 132167 16798 132274
rect 16966 132167 17534 132274
rect 17702 132167 18270 132274
rect 18438 132167 19006 132274
rect 19174 132167 19742 132274
rect 19910 132167 20478 132274
rect 20646 132167 21214 132274
rect 21382 132167 21950 132274
rect 22118 132167 22686 132274
rect 22854 132167 23422 132274
rect 23590 132167 24158 132274
rect 24326 132167 24894 132274
rect 25062 132167 25630 132274
rect 25798 132167 26366 132274
rect 26534 132167 27102 132274
rect 27270 132167 27838 132274
rect 28006 132167 28574 132274
rect 28742 132167 29310 132274
rect 29478 132167 30046 132274
rect 30214 132167 30782 132274
rect 30950 132167 31518 132274
rect 31686 132167 32254 132274
rect 32422 132167 32990 132274
rect 33158 132167 33726 132274
rect 33894 132167 34462 132274
rect 34630 132167 35198 132274
rect 35366 132167 35934 132274
rect 36102 132167 36670 132274
rect 36838 132167 37406 132274
rect 37574 132167 38142 132274
rect 38310 132167 38878 132274
rect 39046 132167 39614 132274
rect 39782 132167 40350 132274
rect 40518 132167 41086 132274
rect 41254 132167 41822 132274
rect 41990 132167 42558 132274
rect 42726 132167 43294 132274
rect 43462 132167 44030 132274
rect 44198 132167 44766 132274
rect 44934 132167 45502 132274
rect 45670 132167 46238 132274
rect 46406 132167 46974 132274
rect 47142 132167 47710 132274
rect 47878 132167 48446 132274
rect 48614 132167 49182 132274
rect 49350 132167 49918 132274
rect 50086 132167 50654 132274
rect 50822 132167 51390 132274
rect 51558 132167 52126 132274
rect 52294 132167 52862 132274
rect 53030 132167 53598 132274
rect 53766 132167 54334 132274
rect 54502 132167 55070 132274
rect 55238 132167 55806 132274
rect 55974 132167 56542 132274
rect 56710 132167 57278 132274
rect 57446 132167 58014 132274
rect 58182 132167 58750 132274
rect 58918 132167 59486 132274
rect 59654 132167 60222 132274
rect 60390 132167 60958 132274
rect 61126 132167 61694 132274
rect 61862 132167 62430 132274
rect 62598 132167 63166 132274
rect 63334 132167 63902 132274
rect 64070 132167 64638 132274
rect 64806 132167 65374 132274
rect 65542 132167 66110 132274
rect 66278 132167 66846 132274
rect 67014 132167 67582 132274
rect 67750 132167 68318 132274
rect 68486 132167 69054 132274
rect 69222 132167 69790 132274
rect 69958 132167 70526 132274
rect 70694 132167 71262 132274
rect 71430 132167 71998 132274
rect 72166 132167 72734 132274
rect 72902 132167 73470 132274
rect 73638 132167 74206 132274
rect 74374 132167 74942 132274
rect 75110 132167 75678 132274
rect 75846 132167 76414 132274
rect 76582 132167 77150 132274
rect 77318 132167 77886 132274
rect 78054 132167 78622 132274
rect 78790 132167 79358 132274
rect 79526 132167 80094 132274
rect 80262 132167 80830 132274
rect 80998 132167 81566 132274
rect 81734 132167 82302 132274
rect 82470 132167 83038 132274
rect 83206 132167 83774 132274
rect 83942 132167 84510 132274
rect 84678 132167 85246 132274
rect 85414 132167 85982 132274
rect 86150 132167 86718 132274
rect 86886 132167 87454 132274
rect 87622 132167 88190 132274
rect 88358 132167 88926 132274
rect 89094 132167 89662 132274
rect 89830 132167 90398 132274
rect 90566 132167 91134 132274
rect 91302 132167 91870 132274
rect 92038 132167 92606 132274
rect 92774 132167 93342 132274
rect 93510 132167 94078 132274
rect 94246 132167 94814 132274
rect 94982 132167 95550 132274
rect 95718 132167 96286 132274
rect 96454 132167 97022 132274
rect 97190 132167 97758 132274
rect 97926 132167 98494 132274
rect 98662 132167 99230 132274
rect 99398 132167 99966 132274
rect 100134 132167 100702 132274
rect 100870 132167 101438 132274
rect 101606 132167 102174 132274
rect 102342 132167 102910 132274
rect 103078 132167 103646 132274
rect 103814 132167 104382 132274
rect 104550 132167 105118 132274
rect 105286 132167 105854 132274
rect 106022 132167 106590 132274
rect 106758 132167 107326 132274
rect 107494 132167 108062 132274
rect 108230 132167 108798 132274
rect 108966 132167 109534 132274
rect 109702 132167 110270 132274
rect 110438 132167 111006 132274
rect 111174 132167 111742 132274
rect 111910 132167 112478 132274
rect 112646 132167 113214 132274
rect 113382 132167 113950 132274
rect 114118 132167 114686 132274
rect 114854 132167 115422 132274
rect 115590 132167 116158 132274
rect 116326 132167 116894 132274
rect 117062 132167 117630 132274
rect 117798 132167 118366 132274
rect 118534 132167 119102 132274
rect 119270 132167 119838 132274
rect 120006 132167 120574 132274
rect 120742 132167 121310 132274
rect 121478 132167 122046 132274
rect 122214 132167 122782 132274
rect 122950 132167 123518 132274
rect 123686 132167 124254 132274
rect 124422 132167 124990 132274
rect 125158 132167 125726 132274
rect 125894 132167 126462 132274
rect 126630 132167 127198 132274
rect 127366 132167 128964 132274
rect 1122 856 128964 132167
rect 1122 439 9990 856
rect 10158 439 10174 856
rect 10342 439 10358 856
rect 10526 439 10542 856
rect 10710 439 10726 856
rect 10894 439 10910 856
rect 11078 439 11094 856
rect 11262 439 11278 856
rect 11446 439 11462 856
rect 11630 439 11646 856
rect 11814 439 11830 856
rect 11998 439 12014 856
rect 12182 439 12198 856
rect 12366 439 12382 856
rect 12550 439 12566 856
rect 12734 439 12750 856
rect 12918 439 12934 856
rect 13102 439 13118 856
rect 13286 439 13302 856
rect 13470 439 13486 856
rect 13654 439 13670 856
rect 13838 439 13854 856
rect 14022 439 14038 856
rect 14206 439 14222 856
rect 14390 439 14406 856
rect 14574 439 14590 856
rect 14758 439 14774 856
rect 14942 439 14958 856
rect 15126 439 15142 856
rect 15310 439 15326 856
rect 15494 439 15510 856
rect 15678 439 15694 856
rect 15862 439 15878 856
rect 16046 439 16062 856
rect 16230 439 16246 856
rect 16414 439 16430 856
rect 16598 439 16614 856
rect 16782 439 16798 856
rect 16966 439 16982 856
rect 17150 439 17166 856
rect 17334 439 17350 856
rect 17518 439 17534 856
rect 17702 439 17718 856
rect 17886 439 17902 856
rect 18070 439 18086 856
rect 18254 439 18270 856
rect 18438 439 18454 856
rect 18622 439 18638 856
rect 18806 439 18822 856
rect 18990 439 19006 856
rect 19174 439 19190 856
rect 19358 439 19374 856
rect 19542 439 19558 856
rect 19726 439 19742 856
rect 19910 439 19926 856
rect 20094 439 20110 856
rect 20278 439 20294 856
rect 20462 439 20478 856
rect 20646 439 20662 856
rect 20830 439 20846 856
rect 21014 439 21030 856
rect 21198 439 21214 856
rect 21382 439 21398 856
rect 21566 439 21582 856
rect 21750 439 21766 856
rect 21934 439 21950 856
rect 22118 439 22134 856
rect 22302 439 22318 856
rect 22486 439 22502 856
rect 22670 439 22686 856
rect 22854 439 22870 856
rect 23038 439 23054 856
rect 23222 439 23238 856
rect 23406 439 23422 856
rect 23590 439 23606 856
rect 23774 439 23790 856
rect 23958 439 23974 856
rect 24142 439 24158 856
rect 24326 439 24342 856
rect 24510 439 24526 856
rect 24694 439 24710 856
rect 24878 439 24894 856
rect 25062 439 25078 856
rect 25246 439 25262 856
rect 25430 439 25446 856
rect 25614 439 25630 856
rect 25798 439 25814 856
rect 25982 439 25998 856
rect 26166 439 26182 856
rect 26350 439 26366 856
rect 26534 439 26550 856
rect 26718 439 26734 856
rect 26902 439 26918 856
rect 27086 439 27102 856
rect 27270 439 27286 856
rect 27454 439 27470 856
rect 27638 439 27654 856
rect 27822 439 27838 856
rect 28006 439 28022 856
rect 28190 439 28206 856
rect 28374 439 28390 856
rect 28558 439 28574 856
rect 28742 439 28758 856
rect 28926 439 28942 856
rect 29110 439 29126 856
rect 29294 439 29310 856
rect 29478 439 29494 856
rect 29662 439 29678 856
rect 29846 439 29862 856
rect 30030 439 30046 856
rect 30214 439 30230 856
rect 30398 439 30414 856
rect 30582 439 30598 856
rect 30766 439 30782 856
rect 30950 439 30966 856
rect 31134 439 31150 856
rect 31318 439 31334 856
rect 31502 439 31518 856
rect 31686 439 31702 856
rect 31870 439 31886 856
rect 32054 439 32070 856
rect 32238 439 32254 856
rect 32422 439 32438 856
rect 32606 439 32622 856
rect 32790 439 32806 856
rect 32974 439 32990 856
rect 33158 439 33174 856
rect 33342 439 33358 856
rect 33526 439 33542 856
rect 33710 439 33726 856
rect 33894 439 33910 856
rect 34078 439 34094 856
rect 34262 439 34278 856
rect 34446 439 34462 856
rect 34630 439 34646 856
rect 34814 439 34830 856
rect 34998 439 35014 856
rect 35182 439 35198 856
rect 35366 439 35382 856
rect 35550 439 35566 856
rect 35734 439 35750 856
rect 35918 439 35934 856
rect 36102 439 36118 856
rect 36286 439 36302 856
rect 36470 439 36486 856
rect 36654 439 36670 856
rect 36838 439 36854 856
rect 37022 439 37038 856
rect 37206 439 37222 856
rect 37390 439 37406 856
rect 37574 439 37590 856
rect 37758 439 37774 856
rect 37942 439 37958 856
rect 38126 439 38142 856
rect 38310 439 38326 856
rect 38494 439 38510 856
rect 38678 439 38694 856
rect 38862 439 38878 856
rect 39046 439 39062 856
rect 39230 439 39246 856
rect 39414 439 39430 856
rect 39598 439 39614 856
rect 39782 439 39798 856
rect 39966 439 39982 856
rect 40150 439 40166 856
rect 40334 439 40350 856
rect 40518 439 40534 856
rect 40702 439 40718 856
rect 40886 439 40902 856
rect 41070 439 41086 856
rect 41254 439 41270 856
rect 41438 439 41454 856
rect 41622 439 41638 856
rect 41806 439 41822 856
rect 41990 439 42006 856
rect 42174 439 42190 856
rect 42358 439 42374 856
rect 42542 439 42558 856
rect 42726 439 42742 856
rect 42910 439 42926 856
rect 43094 439 43110 856
rect 43278 439 43294 856
rect 43462 439 43478 856
rect 43646 439 43662 856
rect 43830 439 43846 856
rect 44014 439 44030 856
rect 44198 439 44214 856
rect 44382 439 44398 856
rect 44566 439 44582 856
rect 44750 439 44766 856
rect 44934 439 44950 856
rect 45118 439 45134 856
rect 45302 439 45318 856
rect 45486 439 45502 856
rect 45670 439 45686 856
rect 45854 439 45870 856
rect 46038 439 46054 856
rect 46222 439 46238 856
rect 46406 439 46422 856
rect 46590 439 46606 856
rect 46774 439 46790 856
rect 46958 439 46974 856
rect 47142 439 47158 856
rect 47326 439 47342 856
rect 47510 439 47526 856
rect 47694 439 47710 856
rect 47878 439 47894 856
rect 48062 439 48078 856
rect 48246 439 48262 856
rect 48430 439 48446 856
rect 48614 439 48630 856
rect 48798 439 48814 856
rect 48982 439 48998 856
rect 49166 439 49182 856
rect 49350 439 49366 856
rect 49534 439 49550 856
rect 49718 439 49734 856
rect 49902 439 49918 856
rect 50086 439 50102 856
rect 50270 439 50286 856
rect 50454 439 50470 856
rect 50638 439 50654 856
rect 50822 439 50838 856
rect 51006 439 51022 856
rect 51190 439 51206 856
rect 51374 439 51390 856
rect 51558 439 51574 856
rect 51742 439 51758 856
rect 51926 439 51942 856
rect 52110 439 52126 856
rect 52294 439 52310 856
rect 52478 439 52494 856
rect 52662 439 52678 856
rect 52846 439 52862 856
rect 53030 439 53046 856
rect 53214 439 53230 856
rect 53398 439 53414 856
rect 53582 439 53598 856
rect 53766 439 53782 856
rect 53950 439 53966 856
rect 54134 439 54150 856
rect 54318 439 54334 856
rect 54502 439 54518 856
rect 54686 439 54702 856
rect 54870 439 54886 856
rect 55054 439 55070 856
rect 55238 439 55254 856
rect 55422 439 55438 856
rect 55606 439 55622 856
rect 55790 439 55806 856
rect 55974 439 55990 856
rect 56158 439 56174 856
rect 56342 439 56358 856
rect 56526 439 56542 856
rect 56710 439 56726 856
rect 56894 439 56910 856
rect 57078 439 57094 856
rect 57262 439 57278 856
rect 57446 439 57462 856
rect 57630 439 57646 856
rect 57814 439 57830 856
rect 57998 439 58014 856
rect 58182 439 58198 856
rect 58366 439 58382 856
rect 58550 439 58566 856
rect 58734 439 58750 856
rect 58918 439 58934 856
rect 59102 439 59118 856
rect 59286 439 59302 856
rect 59470 439 59486 856
rect 59654 439 59670 856
rect 59838 439 59854 856
rect 60022 439 60038 856
rect 60206 439 60222 856
rect 60390 439 60406 856
rect 60574 439 60590 856
rect 60758 439 60774 856
rect 60942 439 60958 856
rect 61126 439 61142 856
rect 61310 439 61326 856
rect 61494 439 61510 856
rect 61678 439 61694 856
rect 61862 439 61878 856
rect 62046 439 62062 856
rect 62230 439 62246 856
rect 62414 439 62430 856
rect 62598 439 62614 856
rect 62782 439 62798 856
rect 62966 439 62982 856
rect 63150 439 63166 856
rect 63334 439 63350 856
rect 63518 439 63534 856
rect 63702 439 63718 856
rect 63886 439 63902 856
rect 64070 439 64086 856
rect 64254 439 64270 856
rect 64438 439 64454 856
rect 64622 439 64638 856
rect 64806 439 64822 856
rect 64990 439 65006 856
rect 65174 439 65190 856
rect 65358 439 65374 856
rect 65542 439 65558 856
rect 65726 439 65742 856
rect 65910 439 65926 856
rect 66094 439 66110 856
rect 66278 439 66294 856
rect 66462 439 66478 856
rect 66646 439 66662 856
rect 66830 439 66846 856
rect 67014 439 67030 856
rect 67198 439 67214 856
rect 67382 439 67398 856
rect 67566 439 67582 856
rect 67750 439 67766 856
rect 67934 439 67950 856
rect 68118 439 68134 856
rect 68302 439 68318 856
rect 68486 439 68502 856
rect 68670 439 68686 856
rect 68854 439 68870 856
rect 69038 439 69054 856
rect 69222 439 69238 856
rect 69406 439 69422 856
rect 69590 439 69606 856
rect 69774 439 69790 856
rect 69958 439 69974 856
rect 70142 439 70158 856
rect 70326 439 70342 856
rect 70510 439 70526 856
rect 70694 439 70710 856
rect 70878 439 70894 856
rect 71062 439 71078 856
rect 71246 439 71262 856
rect 71430 439 71446 856
rect 71614 439 71630 856
rect 71798 439 71814 856
rect 71982 439 71998 856
rect 72166 439 72182 856
rect 72350 439 72366 856
rect 72534 439 72550 856
rect 72718 439 72734 856
rect 72902 439 72918 856
rect 73086 439 73102 856
rect 73270 439 73286 856
rect 73454 439 73470 856
rect 73638 439 73654 856
rect 73822 439 73838 856
rect 74006 439 74022 856
rect 74190 439 74206 856
rect 74374 439 74390 856
rect 74558 439 74574 856
rect 74742 439 74758 856
rect 74926 439 74942 856
rect 75110 439 75126 856
rect 75294 439 75310 856
rect 75478 439 75494 856
rect 75662 439 75678 856
rect 75846 439 75862 856
rect 76030 439 76046 856
rect 76214 439 76230 856
rect 76398 439 76414 856
rect 76582 439 76598 856
rect 76766 439 76782 856
rect 76950 439 76966 856
rect 77134 439 77150 856
rect 77318 439 77334 856
rect 77502 439 77518 856
rect 77686 439 77702 856
rect 77870 439 77886 856
rect 78054 439 78070 856
rect 78238 439 78254 856
rect 78422 439 78438 856
rect 78606 439 78622 856
rect 78790 439 78806 856
rect 78974 439 78990 856
rect 79158 439 79174 856
rect 79342 439 79358 856
rect 79526 439 79542 856
rect 79710 439 79726 856
rect 79894 439 79910 856
rect 80078 439 80094 856
rect 80262 439 80278 856
rect 80446 439 80462 856
rect 80630 439 80646 856
rect 80814 439 80830 856
rect 80998 439 81014 856
rect 81182 439 81198 856
rect 81366 439 81382 856
rect 81550 439 81566 856
rect 81734 439 81750 856
rect 81918 439 81934 856
rect 82102 439 82118 856
rect 82286 439 82302 856
rect 82470 439 82486 856
rect 82654 439 82670 856
rect 82838 439 82854 856
rect 83022 439 83038 856
rect 83206 439 83222 856
rect 83390 439 83406 856
rect 83574 439 83590 856
rect 83758 439 83774 856
rect 83942 439 83958 856
rect 84126 439 84142 856
rect 84310 439 84326 856
rect 84494 439 84510 856
rect 84678 439 84694 856
rect 84862 439 84878 856
rect 85046 439 85062 856
rect 85230 439 85246 856
rect 85414 439 85430 856
rect 85598 439 85614 856
rect 85782 439 85798 856
rect 85966 439 85982 856
rect 86150 439 86166 856
rect 86334 439 86350 856
rect 86518 439 86534 856
rect 86702 439 86718 856
rect 86886 439 86902 856
rect 87070 439 87086 856
rect 87254 439 87270 856
rect 87438 439 87454 856
rect 87622 439 87638 856
rect 87806 439 87822 856
rect 87990 439 88006 856
rect 88174 439 88190 856
rect 88358 439 88374 856
rect 88542 439 88558 856
rect 88726 439 88742 856
rect 88910 439 88926 856
rect 89094 439 89110 856
rect 89278 439 89294 856
rect 89462 439 89478 856
rect 89646 439 89662 856
rect 89830 439 89846 856
rect 90014 439 90030 856
rect 90198 439 90214 856
rect 90382 439 90398 856
rect 90566 439 90582 856
rect 90750 439 90766 856
rect 90934 439 90950 856
rect 91118 439 91134 856
rect 91302 439 91318 856
rect 91486 439 91502 856
rect 91670 439 91686 856
rect 91854 439 91870 856
rect 92038 439 92054 856
rect 92222 439 92238 856
rect 92406 439 92422 856
rect 92590 439 92606 856
rect 92774 439 92790 856
rect 92958 439 92974 856
rect 93142 439 93158 856
rect 93326 439 93342 856
rect 93510 439 93526 856
rect 93694 439 93710 856
rect 93878 439 93894 856
rect 94062 439 94078 856
rect 94246 439 94262 856
rect 94430 439 94446 856
rect 94614 439 94630 856
rect 94798 439 94814 856
rect 94982 439 94998 856
rect 95166 439 95182 856
rect 95350 439 95366 856
rect 95534 439 95550 856
rect 95718 439 95734 856
rect 95902 439 95918 856
rect 96086 439 96102 856
rect 96270 439 96286 856
rect 96454 439 96470 856
rect 96638 439 96654 856
rect 96822 439 96838 856
rect 97006 439 97022 856
rect 97190 439 97206 856
rect 97374 439 97390 856
rect 97558 439 97574 856
rect 97742 439 97758 856
rect 97926 439 97942 856
rect 98110 439 98126 856
rect 98294 439 98310 856
rect 98478 439 98494 856
rect 98662 439 98678 856
rect 98846 439 98862 856
rect 99030 439 99046 856
rect 99214 439 99230 856
rect 99398 439 99414 856
rect 99582 439 99598 856
rect 99766 439 99782 856
rect 99950 439 99966 856
rect 100134 439 100150 856
rect 100318 439 100334 856
rect 100502 439 100518 856
rect 100686 439 100702 856
rect 100870 439 100886 856
rect 101054 439 101070 856
rect 101238 439 101254 856
rect 101422 439 101438 856
rect 101606 439 101622 856
rect 101790 439 101806 856
rect 101974 439 101990 856
rect 102158 439 102174 856
rect 102342 439 102358 856
rect 102526 439 102542 856
rect 102710 439 102726 856
rect 102894 439 102910 856
rect 103078 439 103094 856
rect 103262 439 103278 856
rect 103446 439 103462 856
rect 103630 439 103646 856
rect 103814 439 103830 856
rect 103998 439 104014 856
rect 104182 439 104198 856
rect 104366 439 104382 856
rect 104550 439 104566 856
rect 104734 439 104750 856
rect 104918 439 104934 856
rect 105102 439 105118 856
rect 105286 439 105302 856
rect 105470 439 105486 856
rect 105654 439 105670 856
rect 105838 439 105854 856
rect 106022 439 106038 856
rect 106206 439 106222 856
rect 106390 439 106406 856
rect 106574 439 106590 856
rect 106758 439 106774 856
rect 106942 439 106958 856
rect 107126 439 107142 856
rect 107310 439 107326 856
rect 107494 439 107510 856
rect 107678 439 107694 856
rect 107862 439 107878 856
rect 108046 439 108062 856
rect 108230 439 108246 856
rect 108414 439 108430 856
rect 108598 439 108614 856
rect 108782 439 108798 856
rect 108966 439 108982 856
rect 109150 439 109166 856
rect 109334 439 109350 856
rect 109518 439 109534 856
rect 109702 439 109718 856
rect 109886 439 109902 856
rect 110070 439 110086 856
rect 110254 439 110270 856
rect 110438 439 110454 856
rect 110622 439 110638 856
rect 110806 439 110822 856
rect 110990 439 111006 856
rect 111174 439 111190 856
rect 111358 439 111374 856
rect 111542 439 111558 856
rect 111726 439 111742 856
rect 111910 439 111926 856
rect 112094 439 112110 856
rect 112278 439 112294 856
rect 112462 439 112478 856
rect 112646 439 112662 856
rect 112830 439 112846 856
rect 113014 439 113030 856
rect 113198 439 113214 856
rect 113382 439 113398 856
rect 113566 439 113582 856
rect 113750 439 113766 856
rect 113934 439 113950 856
rect 114118 439 114134 856
rect 114302 439 114318 856
rect 114486 439 114502 856
rect 114670 439 114686 856
rect 114854 439 114870 856
rect 115038 439 115054 856
rect 115222 439 115238 856
rect 115406 439 115422 856
rect 115590 439 115606 856
rect 115774 439 115790 856
rect 115958 439 115974 856
rect 116142 439 116158 856
rect 116326 439 116342 856
rect 116510 439 116526 856
rect 116694 439 116710 856
rect 116878 439 116894 856
rect 117062 439 117078 856
rect 117246 439 117262 856
rect 117430 439 117446 856
rect 117614 439 117630 856
rect 117798 439 117814 856
rect 117982 439 117998 856
rect 118166 439 118182 856
rect 118350 439 118366 856
rect 118534 439 118550 856
rect 118718 439 118734 856
rect 118902 439 118918 856
rect 119086 439 119102 856
rect 119270 439 119286 856
rect 119454 439 119470 856
rect 119638 439 119654 856
rect 119822 439 119838 856
rect 120006 439 120022 856
rect 120190 439 120206 856
rect 120374 439 120390 856
rect 120558 439 120574 856
rect 120742 439 120758 856
rect 120926 439 128964 856
<< obsm3 >>
rect 1117 443 127959 130797
<< metal4 >>
rect 4208 2128 4528 130608
rect 19568 2128 19888 130608
rect 34928 2128 35248 130608
rect 50288 2128 50608 130608
rect 65648 2128 65968 130608
rect 81008 2128 81328 130608
rect 96368 2128 96688 130608
rect 111728 2128 112048 130608
rect 127088 2128 127408 130608
<< obsm4 >>
rect 2819 130688 126901 130797
rect 2819 2048 4128 130688
rect 4608 2048 19488 130688
rect 19968 2048 34848 130688
rect 35328 2048 50208 130688
rect 50688 2048 65568 130688
rect 66048 2048 80928 130688
rect 81408 2048 96288 130688
rect 96768 2048 111648 130688
rect 112128 2048 126901 130688
rect 2819 443 126901 2048
<< labels >>
rlabel metal2 s 5814 132223 5870 133023 6 dram_addr0[0]
port 1 nsew signal output
rlabel metal2 s 8758 132223 8814 133023 6 dram_addr0[1]
port 2 nsew signal output
rlabel metal2 s 11702 132223 11758 133023 6 dram_addr0[2]
port 3 nsew signal output
rlabel metal2 s 14646 132223 14702 133023 6 dram_addr0[3]
port 4 nsew signal output
rlabel metal2 s 17590 132223 17646 133023 6 dram_addr0[4]
port 5 nsew signal output
rlabel metal2 s 19798 132223 19854 133023 6 dram_addr0[5]
port 6 nsew signal output
rlabel metal2 s 22006 132223 22062 133023 6 dram_addr0[6]
port 7 nsew signal output
rlabel metal2 s 24214 132223 24270 133023 6 dram_addr0[7]
port 8 nsew signal output
rlabel metal2 s 26422 132223 26478 133023 6 dram_addr0[8]
port 9 nsew signal output
rlabel metal2 s 3606 132223 3662 133023 6 dram_clk0
port 10 nsew signal output
rlabel metal2 s 4342 132223 4398 133023 6 dram_csb0
port 11 nsew signal output
rlabel metal2 s 6550 132223 6606 133023 6 dram_din0[0]
port 12 nsew signal output
rlabel metal2 s 30102 132223 30158 133023 6 dram_din0[10]
port 13 nsew signal output
rlabel metal2 s 31574 132223 31630 133023 6 dram_din0[11]
port 14 nsew signal output
rlabel metal2 s 33046 132223 33102 133023 6 dram_din0[12]
port 15 nsew signal output
rlabel metal2 s 34518 132223 34574 133023 6 dram_din0[13]
port 16 nsew signal output
rlabel metal2 s 35990 132223 36046 133023 6 dram_din0[14]
port 17 nsew signal output
rlabel metal2 s 37462 132223 37518 133023 6 dram_din0[15]
port 18 nsew signal output
rlabel metal2 s 38934 132223 38990 133023 6 dram_din0[16]
port 19 nsew signal output
rlabel metal2 s 40406 132223 40462 133023 6 dram_din0[17]
port 20 nsew signal output
rlabel metal2 s 41878 132223 41934 133023 6 dram_din0[18]
port 21 nsew signal output
rlabel metal2 s 43350 132223 43406 133023 6 dram_din0[19]
port 22 nsew signal output
rlabel metal2 s 9494 132223 9550 133023 6 dram_din0[1]
port 23 nsew signal output
rlabel metal2 s 44822 132223 44878 133023 6 dram_din0[20]
port 24 nsew signal output
rlabel metal2 s 46294 132223 46350 133023 6 dram_din0[21]
port 25 nsew signal output
rlabel metal2 s 47766 132223 47822 133023 6 dram_din0[22]
port 26 nsew signal output
rlabel metal2 s 49238 132223 49294 133023 6 dram_din0[23]
port 27 nsew signal output
rlabel metal2 s 50710 132223 50766 133023 6 dram_din0[24]
port 28 nsew signal output
rlabel metal2 s 52182 132223 52238 133023 6 dram_din0[25]
port 29 nsew signal output
rlabel metal2 s 53654 132223 53710 133023 6 dram_din0[26]
port 30 nsew signal output
rlabel metal2 s 55126 132223 55182 133023 6 dram_din0[27]
port 31 nsew signal output
rlabel metal2 s 56598 132223 56654 133023 6 dram_din0[28]
port 32 nsew signal output
rlabel metal2 s 58070 132223 58126 133023 6 dram_din0[29]
port 33 nsew signal output
rlabel metal2 s 12438 132223 12494 133023 6 dram_din0[2]
port 34 nsew signal output
rlabel metal2 s 59542 132223 59598 133023 6 dram_din0[30]
port 35 nsew signal output
rlabel metal2 s 61014 132223 61070 133023 6 dram_din0[31]
port 36 nsew signal output
rlabel metal2 s 15382 132223 15438 133023 6 dram_din0[3]
port 37 nsew signal output
rlabel metal2 s 18326 132223 18382 133023 6 dram_din0[4]
port 38 nsew signal output
rlabel metal2 s 20534 132223 20590 133023 6 dram_din0[5]
port 39 nsew signal output
rlabel metal2 s 22742 132223 22798 133023 6 dram_din0[6]
port 40 nsew signal output
rlabel metal2 s 24950 132223 25006 133023 6 dram_din0[7]
port 41 nsew signal output
rlabel metal2 s 27158 132223 27214 133023 6 dram_din0[8]
port 42 nsew signal output
rlabel metal2 s 28630 132223 28686 133023 6 dram_din0[9]
port 43 nsew signal output
rlabel metal2 s 7286 132223 7342 133023 6 dram_dout0[0]
port 44 nsew signal input
rlabel metal2 s 30838 132223 30894 133023 6 dram_dout0[10]
port 45 nsew signal input
rlabel metal2 s 32310 132223 32366 133023 6 dram_dout0[11]
port 46 nsew signal input
rlabel metal2 s 33782 132223 33838 133023 6 dram_dout0[12]
port 47 nsew signal input
rlabel metal2 s 35254 132223 35310 133023 6 dram_dout0[13]
port 48 nsew signal input
rlabel metal2 s 36726 132223 36782 133023 6 dram_dout0[14]
port 49 nsew signal input
rlabel metal2 s 38198 132223 38254 133023 6 dram_dout0[15]
port 50 nsew signal input
rlabel metal2 s 39670 132223 39726 133023 6 dram_dout0[16]
port 51 nsew signal input
rlabel metal2 s 41142 132223 41198 133023 6 dram_dout0[17]
port 52 nsew signal input
rlabel metal2 s 42614 132223 42670 133023 6 dram_dout0[18]
port 53 nsew signal input
rlabel metal2 s 44086 132223 44142 133023 6 dram_dout0[19]
port 54 nsew signal input
rlabel metal2 s 10230 132223 10286 133023 6 dram_dout0[1]
port 55 nsew signal input
rlabel metal2 s 45558 132223 45614 133023 6 dram_dout0[20]
port 56 nsew signal input
rlabel metal2 s 47030 132223 47086 133023 6 dram_dout0[21]
port 57 nsew signal input
rlabel metal2 s 48502 132223 48558 133023 6 dram_dout0[22]
port 58 nsew signal input
rlabel metal2 s 49974 132223 50030 133023 6 dram_dout0[23]
port 59 nsew signal input
rlabel metal2 s 51446 132223 51502 133023 6 dram_dout0[24]
port 60 nsew signal input
rlabel metal2 s 52918 132223 52974 133023 6 dram_dout0[25]
port 61 nsew signal input
rlabel metal2 s 54390 132223 54446 133023 6 dram_dout0[26]
port 62 nsew signal input
rlabel metal2 s 55862 132223 55918 133023 6 dram_dout0[27]
port 63 nsew signal input
rlabel metal2 s 57334 132223 57390 133023 6 dram_dout0[28]
port 64 nsew signal input
rlabel metal2 s 58806 132223 58862 133023 6 dram_dout0[29]
port 65 nsew signal input
rlabel metal2 s 13174 132223 13230 133023 6 dram_dout0[2]
port 66 nsew signal input
rlabel metal2 s 60278 132223 60334 133023 6 dram_dout0[30]
port 67 nsew signal input
rlabel metal2 s 61750 132223 61806 133023 6 dram_dout0[31]
port 68 nsew signal input
rlabel metal2 s 16118 132223 16174 133023 6 dram_dout0[3]
port 69 nsew signal input
rlabel metal2 s 19062 132223 19118 133023 6 dram_dout0[4]
port 70 nsew signal input
rlabel metal2 s 21270 132223 21326 133023 6 dram_dout0[5]
port 71 nsew signal input
rlabel metal2 s 23478 132223 23534 133023 6 dram_dout0[6]
port 72 nsew signal input
rlabel metal2 s 25686 132223 25742 133023 6 dram_dout0[7]
port 73 nsew signal input
rlabel metal2 s 27894 132223 27950 133023 6 dram_dout0[8]
port 74 nsew signal input
rlabel metal2 s 29366 132223 29422 133023 6 dram_dout0[9]
port 75 nsew signal input
rlabel metal2 s 5078 132223 5134 133023 6 dram_web0
port 76 nsew signal output
rlabel metal2 s 8022 132223 8078 133023 6 dram_wmask0[0]
port 77 nsew signal output
rlabel metal2 s 10966 132223 11022 133023 6 dram_wmask0[1]
port 78 nsew signal output
rlabel metal2 s 13910 132223 13966 133023 6 dram_wmask0[2]
port 79 nsew signal output
rlabel metal2 s 16854 132223 16910 133023 6 dram_wmask0[3]
port 80 nsew signal output
rlabel metal2 s 64694 132223 64750 133023 6 gpio_in[0]
port 81 nsew signal input
rlabel metal2 s 86774 132223 86830 133023 6 gpio_in[10]
port 82 nsew signal input
rlabel metal2 s 88982 132223 89038 133023 6 gpio_in[11]
port 83 nsew signal input
rlabel metal2 s 91190 132223 91246 133023 6 gpio_in[12]
port 84 nsew signal input
rlabel metal2 s 93398 132223 93454 133023 6 gpio_in[13]
port 85 nsew signal input
rlabel metal2 s 95606 132223 95662 133023 6 gpio_in[14]
port 86 nsew signal input
rlabel metal2 s 97814 132223 97870 133023 6 gpio_in[15]
port 87 nsew signal input
rlabel metal2 s 100022 132223 100078 133023 6 gpio_in[16]
port 88 nsew signal input
rlabel metal2 s 102230 132223 102286 133023 6 gpio_in[17]
port 89 nsew signal input
rlabel metal2 s 104438 132223 104494 133023 6 gpio_in[18]
port 90 nsew signal input
rlabel metal2 s 106646 132223 106702 133023 6 gpio_in[19]
port 91 nsew signal input
rlabel metal2 s 66902 132223 66958 133023 6 gpio_in[1]
port 92 nsew signal input
rlabel metal2 s 108854 132223 108910 133023 6 gpio_in[20]
port 93 nsew signal input
rlabel metal2 s 111062 132223 111118 133023 6 gpio_in[21]
port 94 nsew signal input
rlabel metal2 s 113270 132223 113326 133023 6 gpio_in[22]
port 95 nsew signal input
rlabel metal2 s 115478 132223 115534 133023 6 gpio_in[23]
port 96 nsew signal input
rlabel metal2 s 69110 132223 69166 133023 6 gpio_in[2]
port 97 nsew signal input
rlabel metal2 s 71318 132223 71374 133023 6 gpio_in[3]
port 98 nsew signal input
rlabel metal2 s 73526 132223 73582 133023 6 gpio_in[4]
port 99 nsew signal input
rlabel metal2 s 75734 132223 75790 133023 6 gpio_in[5]
port 100 nsew signal input
rlabel metal2 s 77942 132223 77998 133023 6 gpio_in[6]
port 101 nsew signal input
rlabel metal2 s 80150 132223 80206 133023 6 gpio_in[7]
port 102 nsew signal input
rlabel metal2 s 82358 132223 82414 133023 6 gpio_in[8]
port 103 nsew signal input
rlabel metal2 s 84566 132223 84622 133023 6 gpio_in[9]
port 104 nsew signal input
rlabel metal2 s 65430 132223 65486 133023 6 gpio_oeb[0]
port 105 nsew signal output
rlabel metal2 s 87510 132223 87566 133023 6 gpio_oeb[10]
port 106 nsew signal output
rlabel metal2 s 89718 132223 89774 133023 6 gpio_oeb[11]
port 107 nsew signal output
rlabel metal2 s 91926 132223 91982 133023 6 gpio_oeb[12]
port 108 nsew signal output
rlabel metal2 s 94134 132223 94190 133023 6 gpio_oeb[13]
port 109 nsew signal output
rlabel metal2 s 96342 132223 96398 133023 6 gpio_oeb[14]
port 110 nsew signal output
rlabel metal2 s 98550 132223 98606 133023 6 gpio_oeb[15]
port 111 nsew signal output
rlabel metal2 s 100758 132223 100814 133023 6 gpio_oeb[16]
port 112 nsew signal output
rlabel metal2 s 102966 132223 103022 133023 6 gpio_oeb[17]
port 113 nsew signal output
rlabel metal2 s 105174 132223 105230 133023 6 gpio_oeb[18]
port 114 nsew signal output
rlabel metal2 s 107382 132223 107438 133023 6 gpio_oeb[19]
port 115 nsew signal output
rlabel metal2 s 67638 132223 67694 133023 6 gpio_oeb[1]
port 116 nsew signal output
rlabel metal2 s 109590 132223 109646 133023 6 gpio_oeb[20]
port 117 nsew signal output
rlabel metal2 s 111798 132223 111854 133023 6 gpio_oeb[21]
port 118 nsew signal output
rlabel metal2 s 114006 132223 114062 133023 6 gpio_oeb[22]
port 119 nsew signal output
rlabel metal2 s 116214 132223 116270 133023 6 gpio_oeb[23]
port 120 nsew signal output
rlabel metal2 s 117686 132223 117742 133023 6 gpio_oeb[24]
port 121 nsew signal output
rlabel metal2 s 118422 132223 118478 133023 6 gpio_oeb[25]
port 122 nsew signal output
rlabel metal2 s 119158 132223 119214 133023 6 gpio_oeb[26]
port 123 nsew signal output
rlabel metal2 s 119894 132223 119950 133023 6 gpio_oeb[27]
port 124 nsew signal output
rlabel metal2 s 120630 132223 120686 133023 6 gpio_oeb[28]
port 125 nsew signal output
rlabel metal2 s 121366 132223 121422 133023 6 gpio_oeb[29]
port 126 nsew signal output
rlabel metal2 s 69846 132223 69902 133023 6 gpio_oeb[2]
port 127 nsew signal output
rlabel metal2 s 122102 132223 122158 133023 6 gpio_oeb[30]
port 128 nsew signal output
rlabel metal2 s 122838 132223 122894 133023 6 gpio_oeb[31]
port 129 nsew signal output
rlabel metal2 s 123574 132223 123630 133023 6 gpio_oeb[32]
port 130 nsew signal output
rlabel metal2 s 124310 132223 124366 133023 6 gpio_oeb[33]
port 131 nsew signal output
rlabel metal2 s 125046 132223 125102 133023 6 gpio_oeb[34]
port 132 nsew signal output
rlabel metal2 s 125782 132223 125838 133023 6 gpio_oeb[35]
port 133 nsew signal output
rlabel metal2 s 126518 132223 126574 133023 6 gpio_oeb[36]
port 134 nsew signal output
rlabel metal2 s 127254 132223 127310 133023 6 gpio_oeb[37]
port 135 nsew signal output
rlabel metal2 s 72054 132223 72110 133023 6 gpio_oeb[3]
port 136 nsew signal output
rlabel metal2 s 74262 132223 74318 133023 6 gpio_oeb[4]
port 137 nsew signal output
rlabel metal2 s 76470 132223 76526 133023 6 gpio_oeb[5]
port 138 nsew signal output
rlabel metal2 s 78678 132223 78734 133023 6 gpio_oeb[6]
port 139 nsew signal output
rlabel metal2 s 80886 132223 80942 133023 6 gpio_oeb[7]
port 140 nsew signal output
rlabel metal2 s 83094 132223 83150 133023 6 gpio_oeb[8]
port 141 nsew signal output
rlabel metal2 s 85302 132223 85358 133023 6 gpio_oeb[9]
port 142 nsew signal output
rlabel metal2 s 66166 132223 66222 133023 6 gpio_out[0]
port 143 nsew signal output
rlabel metal2 s 88246 132223 88302 133023 6 gpio_out[10]
port 144 nsew signal output
rlabel metal2 s 90454 132223 90510 133023 6 gpio_out[11]
port 145 nsew signal output
rlabel metal2 s 92662 132223 92718 133023 6 gpio_out[12]
port 146 nsew signal output
rlabel metal2 s 94870 132223 94926 133023 6 gpio_out[13]
port 147 nsew signal output
rlabel metal2 s 97078 132223 97134 133023 6 gpio_out[14]
port 148 nsew signal output
rlabel metal2 s 99286 132223 99342 133023 6 gpio_out[15]
port 149 nsew signal output
rlabel metal2 s 101494 132223 101550 133023 6 gpio_out[16]
port 150 nsew signal output
rlabel metal2 s 103702 132223 103758 133023 6 gpio_out[17]
port 151 nsew signal output
rlabel metal2 s 105910 132223 105966 133023 6 gpio_out[18]
port 152 nsew signal output
rlabel metal2 s 108118 132223 108174 133023 6 gpio_out[19]
port 153 nsew signal output
rlabel metal2 s 68374 132223 68430 133023 6 gpio_out[1]
port 154 nsew signal output
rlabel metal2 s 110326 132223 110382 133023 6 gpio_out[20]
port 155 nsew signal output
rlabel metal2 s 112534 132223 112590 133023 6 gpio_out[21]
port 156 nsew signal output
rlabel metal2 s 114742 132223 114798 133023 6 gpio_out[22]
port 157 nsew signal output
rlabel metal2 s 116950 132223 117006 133023 6 gpio_out[23]
port 158 nsew signal output
rlabel metal2 s 70582 132223 70638 133023 6 gpio_out[2]
port 159 nsew signal output
rlabel metal2 s 72790 132223 72846 133023 6 gpio_out[3]
port 160 nsew signal output
rlabel metal2 s 74998 132223 75054 133023 6 gpio_out[4]
port 161 nsew signal output
rlabel metal2 s 77206 132223 77262 133023 6 gpio_out[5]
port 162 nsew signal output
rlabel metal2 s 79414 132223 79470 133023 6 gpio_out[6]
port 163 nsew signal output
rlabel metal2 s 81622 132223 81678 133023 6 gpio_out[7]
port 164 nsew signal output
rlabel metal2 s 83830 132223 83886 133023 6 gpio_out[8]
port 165 nsew signal output
rlabel metal2 s 86038 132223 86094 133023 6 gpio_out[9]
port 166 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 iram_addr0[0]
port 167 nsew signal output
rlabel metal2 s 101862 0 101918 800 6 iram_addr0[1]
port 168 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 iram_addr0[2]
port 169 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 iram_addr0[3]
port 170 nsew signal output
rlabel metal2 s 104622 0 104678 800 6 iram_addr0[4]
port 171 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 iram_addr0[5]
port 172 nsew signal output
rlabel metal2 s 106094 0 106150 800 6 iram_addr0[6]
port 173 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 iram_addr0[7]
port 174 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 iram_addr0[8]
port 175 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 iram_clk0
port 176 nsew signal output
rlabel metal2 s 100390 0 100446 800 6 iram_csb0_A
port 177 nsew signal output
rlabel metal2 s 100574 0 100630 800 6 iram_csb0_B
port 178 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 iram_din0[0]
port 179 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 iram_din0[10]
port 180 nsew signal output
rlabel metal2 s 109406 0 109462 800 6 iram_din0[11]
port 181 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 iram_din0[12]
port 182 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 iram_din0[13]
port 183 nsew signal output
rlabel metal2 s 111062 0 111118 800 6 iram_din0[14]
port 184 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 iram_din0[15]
port 185 nsew signal output
rlabel metal2 s 112166 0 112222 800 6 iram_din0[16]
port 186 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 iram_din0[17]
port 187 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 iram_din0[18]
port 188 nsew signal output
rlabel metal2 s 113822 0 113878 800 6 iram_din0[19]
port 189 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 iram_din0[1]
port 190 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 iram_din0[20]
port 191 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 iram_din0[21]
port 192 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 iram_din0[22]
port 193 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 iram_din0[23]
port 194 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 iram_din0[24]
port 195 nsew signal output
rlabel metal2 s 117134 0 117190 800 6 iram_din0[25]
port 196 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 iram_din0[26]
port 197 nsew signal output
rlabel metal2 s 118238 0 118294 800 6 iram_din0[27]
port 198 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 iram_din0[28]
port 199 nsew signal output
rlabel metal2 s 119342 0 119398 800 6 iram_din0[29]
port 200 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 iram_din0[2]
port 201 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 iram_din0[30]
port 202 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 iram_din0[31]
port 203 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 iram_din0[3]
port 204 nsew signal output
rlabel metal2 s 104806 0 104862 800 6 iram_din0[4]
port 205 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 iram_din0[5]
port 206 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 iram_din0[6]
port 207 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 iram_din0[7]
port 208 nsew signal output
rlabel metal2 s 107750 0 107806 800 6 iram_din0[8]
port 209 nsew signal output
rlabel metal2 s 108302 0 108358 800 6 iram_din0[9]
port 210 nsew signal output
rlabel metal2 s 101310 0 101366 800 6 iram_dout0_A[0]
port 211 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 iram_dout0_A[10]
port 212 nsew signal input
rlabel metal2 s 109590 0 109646 800 6 iram_dout0_A[11]
port 213 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 iram_dout0_A[12]
port 214 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 iram_dout0_A[13]
port 215 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 iram_dout0_A[14]
port 216 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 iram_dout0_A[15]
port 217 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 iram_dout0_A[16]
port 218 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 iram_dout0_A[17]
port 219 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 iram_dout0_A[18]
port 220 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 iram_dout0_A[19]
port 221 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 iram_dout0_A[1]
port 222 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 iram_dout0_A[20]
port 223 nsew signal input
rlabel metal2 s 115110 0 115166 800 6 iram_dout0_A[21]
port 224 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 iram_dout0_A[22]
port 225 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 iram_dout0_A[23]
port 226 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 iram_dout0_A[24]
port 227 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 iram_dout0_A[25]
port 228 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 iram_dout0_A[26]
port 229 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 iram_dout0_A[27]
port 230 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 iram_dout0_A[28]
port 231 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 iram_dout0_A[29]
port 232 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 iram_dout0_A[2]
port 233 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 iram_dout0_A[30]
port 234 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 iram_dout0_A[31]
port 235 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 iram_dout0_A[3]
port 236 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 iram_dout0_A[4]
port 237 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 iram_dout0_A[5]
port 238 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 iram_dout0_A[6]
port 239 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 iram_dout0_A[7]
port 240 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 iram_dout0_A[8]
port 241 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 iram_dout0_A[9]
port 242 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 iram_dout0_B[0]
port 243 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 iram_dout0_B[10]
port 244 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 iram_dout0_B[11]
port 245 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 iram_dout0_B[12]
port 246 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 iram_dout0_B[13]
port 247 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 iram_dout0_B[14]
port 248 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 iram_dout0_B[15]
port 249 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 iram_dout0_B[16]
port 250 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 iram_dout0_B[17]
port 251 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 iram_dout0_B[18]
port 252 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 iram_dout0_B[19]
port 253 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 iram_dout0_B[1]
port 254 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 iram_dout0_B[20]
port 255 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 iram_dout0_B[21]
port 256 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 iram_dout0_B[22]
port 257 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 iram_dout0_B[23]
port 258 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 iram_dout0_B[24]
port 259 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 iram_dout0_B[25]
port 260 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 iram_dout0_B[26]
port 261 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 iram_dout0_B[27]
port 262 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 iram_dout0_B[28]
port 263 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 iram_dout0_B[29]
port 264 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 iram_dout0_B[2]
port 265 nsew signal input
rlabel metal2 s 120262 0 120318 800 6 iram_dout0_B[30]
port 266 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 iram_dout0_B[31]
port 267 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 iram_dout0_B[3]
port 268 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 iram_dout0_B[4]
port 269 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 iram_dout0_B[5]
port 270 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 iram_dout0_B[6]
port 271 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 iram_dout0_B[7]
port 272 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 iram_dout0_B[8]
port 273 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 iram_dout0_B[9]
port 274 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 iram_web0
port 275 nsew signal output
rlabel metal2 s 101678 0 101734 800 6 iram_wmask0[0]
port 276 nsew signal output
rlabel metal2 s 102598 0 102654 800 6 iram_wmask0[1]
port 277 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 iram_wmask0[2]
port 278 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 iram_wmask0[3]
port 279 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 la_data_in[0]
port 280 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_data_in[100]
port 281 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[101]
port 282 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_data_in[102]
port 283 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[103]
port 284 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[104]
port 285 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[105]
port 286 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_data_in[106]
port 287 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[107]
port 288 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[108]
port 289 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[109]
port 290 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_data_in[10]
port 291 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[110]
port 292 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_data_in[111]
port 293 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_data_in[112]
port 294 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[113]
port 295 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_data_in[114]
port 296 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[115]
port 297 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[116]
port 298 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_data_in[117]
port 299 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_data_in[118]
port 300 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[119]
port 301 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_data_in[11]
port 302 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[120]
port 303 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_data_in[121]
port 304 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_data_in[122]
port 305 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[123]
port 306 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_data_in[124]
port 307 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[125]
port 308 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_data_in[126]
port 309 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_data_in[127]
port 310 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 la_data_in[12]
port 311 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_data_in[13]
port 312 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_data_in[14]
port 313 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_data_in[15]
port 314 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_data_in[16]
port 315 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_data_in[17]
port 316 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_data_in[18]
port 317 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[19]
port 318 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 la_data_in[1]
port 319 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_data_in[20]
port 320 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[21]
port 321 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[22]
port 322 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[23]
port 323 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_data_in[24]
port 324 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_data_in[25]
port 325 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in[26]
port 326 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[27]
port 327 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_data_in[28]
port 328 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_data_in[29]
port 329 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 la_data_in[2]
port 330 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_data_in[30]
port 331 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_data_in[31]
port 332 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_data_in[32]
port 333 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[33]
port 334 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_data_in[34]
port 335 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_data_in[35]
port 336 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_data_in[36]
port 337 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_data_in[37]
port 338 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_data_in[38]
port 339 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_data_in[39]
port 340 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_data_in[3]
port 341 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_data_in[40]
port 342 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_data_in[41]
port 343 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_data_in[42]
port 344 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[43]
port 345 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_data_in[44]
port 346 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_data_in[45]
port 347 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[46]
port 348 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_data_in[47]
port 349 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[48]
port 350 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_data_in[49]
port 351 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_data_in[4]
port 352 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_data_in[50]
port 353 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[51]
port 354 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_data_in[52]
port 355 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[53]
port 356 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_data_in[54]
port 357 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_data_in[55]
port 358 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[56]
port 359 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 la_data_in[57]
port 360 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_data_in[58]
port 361 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_data_in[59]
port 362 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_data_in[5]
port 363 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_data_in[60]
port 364 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_data_in[61]
port 365 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 la_data_in[62]
port 366 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_data_in[63]
port 367 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_data_in[64]
port 368 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[65]
port 369 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[66]
port 370 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_data_in[67]
port 371 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_data_in[68]
port 372 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[69]
port 373 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la_data_in[6]
port 374 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_data_in[70]
port 375 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 la_data_in[71]
port 376 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_data_in[72]
port 377 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_data_in[73]
port 378 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[74]
port 379 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[75]
port 380 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_data_in[76]
port 381 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[77]
port 382 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_data_in[78]
port 383 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[79]
port 384 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 la_data_in[7]
port 385 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[80]
port 386 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_data_in[81]
port 387 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_data_in[82]
port 388 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_data_in[83]
port 389 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[84]
port 390 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[85]
port 391 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_data_in[86]
port 392 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[87]
port 393 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_data_in[88]
port 394 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_data_in[89]
port 395 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_data_in[8]
port 396 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_data_in[90]
port 397 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_data_in[91]
port 398 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_data_in[92]
port 399 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_data_in[93]
port 400 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_data_in[94]
port 401 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_data_in[95]
port 402 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_data_in[96]
port 403 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[97]
port 404 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[98]
port 405 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[99]
port 406 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in[9]
port 407 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_data_out[0]
port 408 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 la_data_out[100]
port 409 nsew signal output
rlabel metal2 s 85486 0 85542 800 6 la_data_out[101]
port 410 nsew signal output
rlabel metal2 s 86038 0 86094 800 6 la_data_out[102]
port 411 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 la_data_out[103]
port 412 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 la_data_out[104]
port 413 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[105]
port 414 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[106]
port 415 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[107]
port 416 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[108]
port 417 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[109]
port 418 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 la_data_out[10]
port 419 nsew signal output
rlabel metal2 s 90454 0 90510 800 6 la_data_out[110]
port 420 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[111]
port 421 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 la_data_out[112]
port 422 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 la_data_out[113]
port 423 nsew signal output
rlabel metal2 s 92662 0 92718 800 6 la_data_out[114]
port 424 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 la_data_out[115]
port 425 nsew signal output
rlabel metal2 s 93766 0 93822 800 6 la_data_out[116]
port 426 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[117]
port 427 nsew signal output
rlabel metal2 s 94870 0 94926 800 6 la_data_out[118]
port 428 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 la_data_out[119]
port 429 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 la_data_out[11]
port 430 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 la_data_out[120]
port 431 nsew signal output
rlabel metal2 s 96526 0 96582 800 6 la_data_out[121]
port 432 nsew signal output
rlabel metal2 s 97078 0 97134 800 6 la_data_out[122]
port 433 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 la_data_out[123]
port 434 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 la_data_out[124]
port 435 nsew signal output
rlabel metal2 s 98734 0 98790 800 6 la_data_out[125]
port 436 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 la_data_out[126]
port 437 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 la_data_out[127]
port 438 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[12]
port 439 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 la_data_out[13]
port 440 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 la_data_out[14]
port 441 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 la_data_out[15]
port 442 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 la_data_out[16]
port 443 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 la_data_out[17]
port 444 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[18]
port 445 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 la_data_out[19]
port 446 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 la_data_out[1]
port 447 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 la_data_out[20]
port 448 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 la_data_out[21]
port 449 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[22]
port 450 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 la_data_out[23]
port 451 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 la_data_out[24]
port 452 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[25]
port 453 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 la_data_out[26]
port 454 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 la_data_out[27]
port 455 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 la_data_out[28]
port 456 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 la_data_out[29]
port 457 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 la_data_out[2]
port 458 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 la_data_out[30]
port 459 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[31]
port 460 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[32]
port 461 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 la_data_out[33]
port 462 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 la_data_out[34]
port 463 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 la_data_out[35]
port 464 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 la_data_out[36]
port 465 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 la_data_out[37]
port 466 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 la_data_out[38]
port 467 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 la_data_out[39]
port 468 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 la_data_out[3]
port 469 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 la_data_out[40]
port 470 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 la_data_out[41]
port 471 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 la_data_out[42]
port 472 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 la_data_out[43]
port 473 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[44]
port 474 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 la_data_out[45]
port 475 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 la_data_out[46]
port 476 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 la_data_out[47]
port 477 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la_data_out[48]
port 478 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 la_data_out[49]
port 479 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 la_data_out[4]
port 480 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 la_data_out[50]
port 481 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[51]
port 482 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 la_data_out[52]
port 483 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[53]
port 484 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 la_data_out[54]
port 485 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 la_data_out[55]
port 486 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 la_data_out[56]
port 487 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 la_data_out[57]
port 488 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la_data_out[58]
port 489 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 la_data_out[59]
port 490 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 la_data_out[5]
port 491 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 la_data_out[60]
port 492 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 la_data_out[61]
port 493 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 la_data_out[62]
port 494 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 la_data_out[63]
port 495 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[64]
port 496 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[65]
port 497 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 la_data_out[66]
port 498 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 la_data_out[67]
port 499 nsew signal output
rlabel metal2 s 67270 0 67326 800 6 la_data_out[68]
port 500 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 la_data_out[69]
port 501 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 la_data_out[6]
port 502 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 la_data_out[70]
port 503 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[71]
port 504 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 la_data_out[72]
port 505 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 la_data_out[73]
port 506 nsew signal output
rlabel metal2 s 70582 0 70638 800 6 la_data_out[74]
port 507 nsew signal output
rlabel metal2 s 71134 0 71190 800 6 la_data_out[75]
port 508 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 la_data_out[76]
port 509 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 la_data_out[77]
port 510 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[78]
port 511 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 la_data_out[79]
port 512 nsew signal output
rlabel metal2 s 33598 0 33654 800 6 la_data_out[7]
port 513 nsew signal output
rlabel metal2 s 73894 0 73950 800 6 la_data_out[80]
port 514 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[81]
port 515 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 la_data_out[82]
port 516 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 la_data_out[83]
port 517 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 la_data_out[84]
port 518 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[85]
port 519 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 la_data_out[86]
port 520 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[87]
port 521 nsew signal output
rlabel metal2 s 78310 0 78366 800 6 la_data_out[88]
port 522 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 la_data_out[89]
port 523 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 la_data_out[8]
port 524 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[90]
port 525 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 la_data_out[91]
port 526 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 la_data_out[92]
port 527 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 la_data_out[93]
port 528 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 la_data_out[94]
port 529 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 la_data_out[95]
port 530 nsew signal output
rlabel metal2 s 82726 0 82782 800 6 la_data_out[96]
port 531 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 la_data_out[97]
port 532 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 la_data_out[98]
port 533 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 la_data_out[99]
port 534 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 la_data_out[9]
port 535 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 la_oenb[0]
port 536 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_oenb[100]
port 537 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_oenb[101]
port 538 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_oenb[102]
port 539 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_oenb[103]
port 540 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_oenb[104]
port 541 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_oenb[105]
port 542 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[106]
port 543 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_oenb[107]
port 544 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 la_oenb[108]
port 545 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_oenb[109]
port 546 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_oenb[10]
port 547 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_oenb[110]
port 548 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_oenb[111]
port 549 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_oenb[112]
port 550 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_oenb[113]
port 551 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_oenb[114]
port 552 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_oenb[115]
port 553 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_oenb[116]
port 554 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_oenb[117]
port 555 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_oenb[118]
port 556 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_oenb[119]
port 557 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 la_oenb[11]
port 558 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_oenb[120]
port 559 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_oenb[121]
port 560 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_oenb[122]
port 561 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_oenb[123]
port 562 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_oenb[124]
port 563 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_oenb[125]
port 564 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_oenb[126]
port 565 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_oenb[127]
port 566 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[12]
port 567 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_oenb[13]
port 568 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 la_oenb[14]
port 569 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 la_oenb[15]
port 570 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_oenb[16]
port 571 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_oenb[17]
port 572 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_oenb[18]
port 573 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_oenb[19]
port 574 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_oenb[1]
port 575 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_oenb[20]
port 576 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_oenb[21]
port 577 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[22]
port 578 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_oenb[23]
port 579 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_oenb[24]
port 580 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_oenb[25]
port 581 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_oenb[26]
port 582 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_oenb[27]
port 583 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_oenb[28]
port 584 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_oenb[29]
port 585 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 la_oenb[2]
port 586 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_oenb[30]
port 587 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_oenb[31]
port 588 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[32]
port 589 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_oenb[33]
port 590 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_oenb[34]
port 591 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_oenb[35]
port 592 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_oenb[36]
port 593 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_oenb[37]
port 594 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_oenb[38]
port 595 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_oenb[39]
port 596 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_oenb[3]
port 597 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_oenb[40]
port 598 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_oenb[41]
port 599 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_oenb[42]
port 600 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oenb[43]
port 601 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_oenb[44]
port 602 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_oenb[45]
port 603 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_oenb[46]
port 604 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_oenb[47]
port 605 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_oenb[48]
port 606 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_oenb[49]
port 607 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 la_oenb[4]
port 608 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oenb[50]
port 609 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_oenb[51]
port 610 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 la_oenb[52]
port 611 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_oenb[53]
port 612 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_oenb[54]
port 613 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[55]
port 614 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_oenb[56]
port 615 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_oenb[57]
port 616 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_oenb[58]
port 617 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_oenb[59]
port 618 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 la_oenb[5]
port 619 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_oenb[60]
port 620 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_oenb[61]
port 621 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_oenb[62]
port 622 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_oenb[63]
port 623 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_oenb[64]
port 624 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[65]
port 625 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_oenb[66]
port 626 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_oenb[67]
port 627 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_oenb[68]
port 628 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_oenb[69]
port 629 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_oenb[6]
port 630 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_oenb[70]
port 631 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 la_oenb[71]
port 632 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_oenb[72]
port 633 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[73]
port 634 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_oenb[74]
port 635 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_oenb[75]
port 636 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_oenb[76]
port 637 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_oenb[77]
port 638 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_oenb[78]
port 639 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oenb[79]
port 640 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 la_oenb[7]
port 641 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[80]
port 642 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oenb[81]
port 643 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_oenb[82]
port 644 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_oenb[83]
port 645 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_oenb[84]
port 646 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 la_oenb[85]
port 647 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_oenb[86]
port 648 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_oenb[87]
port 649 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_oenb[88]
port 650 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_oenb[89]
port 651 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_oenb[8]
port 652 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_oenb[90]
port 653 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_oenb[91]
port 654 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_oenb[92]
port 655 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_oenb[93]
port 656 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[94]
port 657 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[95]
port 658 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 la_oenb[96]
port 659 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[97]
port 660 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oenb[98]
port 661 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_oenb[99]
port 662 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_oenb[9]
port 663 nsew signal input
rlabel metal2 s 62486 132223 62542 133023 6 user_irq[0]
port 664 nsew signal output
rlabel metal2 s 63222 132223 63278 133023 6 user_irq[1]
port 665 nsew signal output
rlabel metal2 s 63958 132223 64014 133023 6 user_irq[2]
port 666 nsew signal output
rlabel metal4 s 4208 2128 4528 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 130608 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 130608 6 vssd1
port 668 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 130608 6 vssd1
port 668 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 130608 6 vssd1
port 668 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 130608 6 vssd1
port 668 nsew ground bidirectional
rlabel metal2 s 10046 0 10102 800 6 wb_clk_i
port 669 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wb_rst_i
port 670 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_ack_o
port 671 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 wbs_adr_i[0]
port 672 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[10]
port 673 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[11]
port 674 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_adr_i[12]
port 675 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[13]
port 676 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_adr_i[14]
port 677 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[15]
port 678 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_adr_i[16]
port 679 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_adr_i[17]
port 680 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_adr_i[18]
port 681 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_adr_i[19]
port 682 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[1]
port 683 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_adr_i[20]
port 684 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_adr_i[21]
port 685 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_adr_i[22]
port 686 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[23]
port 687 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_adr_i[24]
port 688 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_adr_i[25]
port 689 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[26]
port 690 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_adr_i[27]
port 691 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_adr_i[28]
port 692 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_adr_i[29]
port 693 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_adr_i[2]
port 694 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 wbs_adr_i[30]
port 695 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_adr_i[31]
port 696 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[3]
port 697 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_adr_i[4]
port 698 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[5]
port 699 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[6]
port 700 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_adr_i[7]
port 701 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_adr_i[8]
port 702 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_adr_i[9]
port 703 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_cyc_i
port 704 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_i[0]
port 705 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_i[10]
port 706 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[11]
port 707 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[12]
port 708 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[13]
port 709 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_i[14]
port 710 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_i[15]
port 711 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_i[16]
port 712 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[17]
port 713 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_i[18]
port 714 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_i[19]
port 715 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_i[1]
port 716 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_i[20]
port 717 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_i[21]
port 718 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_i[22]
port 719 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_dat_i[23]
port 720 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[24]
port 721 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_i[25]
port 722 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_i[26]
port 723 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_i[27]
port 724 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_i[28]
port 725 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_i[29]
port 726 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_i[2]
port 727 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_i[30]
port 728 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_i[31]
port 729 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_i[3]
port 730 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_i[4]
port 731 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[5]
port 732 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_i[6]
port 733 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_i[7]
port 734 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_i[8]
port 735 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_i[9]
port 736 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_o[0]
port 737 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_o[10]
port 738 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_o[11]
port 739 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[12]
port 740 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_o[13]
port 741 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_o[14]
port 742 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_o[15]
port 743 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_o[16]
port 744 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[17]
port 745 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_o[18]
port 746 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_o[19]
port 747 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_o[1]
port 748 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_o[20]
port 749 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_o[21]
port 750 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_o[22]
port 751 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_o[23]
port 752 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_o[24]
port 753 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_o[25]
port 754 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_o[26]
port 755 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_o[27]
port 756 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_o[28]
port 757 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_o[29]
port 758 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_o[2]
port 759 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_o[30]
port 760 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 wbs_dat_o[31]
port 761 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_o[3]
port 762 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[4]
port 763 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_o[5]
port 764 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_o[6]
port 765 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[7]
port 766 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_o[8]
port 767 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[9]
port 768 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_sel_i[0]
port 769 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_sel_i[1]
port 770 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_sel_i[2]
port 771 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_sel_i[3]
port 772 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_stb_i
port 773 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_we_i
port 774 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 130879 133023
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 43776006
string GDS_FILE /home/jure/Projekti/rvj1-caravel-soc-mpw7/openlane/rvj1_caravel_soc/runs/22_08_08_15_19/results/signoff/rvj1_caravel_soc.magic.gds
string GDS_START 1114732
<< end >>

