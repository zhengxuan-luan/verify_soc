magic
tech sky130A
magscale 1 2
timestamp 1659992954
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 348786 700544 348792 700596
rect 348844 700584 348850 700596
rect 357710 700584 357716 700596
rect 348844 700556 357716 700584
rect 348844 700544 348850 700556
rect 357710 700544 357716 700556
rect 357768 700544 357774 700596
rect 332502 700476 332508 700528
rect 332560 700516 332566 700528
rect 358814 700516 358820 700528
rect 332560 700488 358820 700516
rect 332560 700476 332566 700488
rect 358814 700476 358820 700488
rect 358872 700476 358878 700528
rect 300118 700408 300124 700460
rect 300176 700448 300182 700460
rect 357618 700448 357624 700460
rect 300176 700420 357624 700448
rect 300176 700408 300182 700420
rect 357618 700408 357624 700420
rect 357676 700408 357682 700460
rect 283834 700340 283840 700392
rect 283892 700380 283898 700392
rect 357526 700380 357532 700392
rect 283892 700352 357532 700380
rect 283892 700340 283898 700352
rect 357526 700340 357532 700352
rect 357584 700340 357590 700392
rect 217962 700272 217968 700324
rect 218020 700312 218026 700324
rect 235166 700312 235172 700324
rect 218020 700284 235172 700312
rect 218020 700272 218026 700284
rect 235166 700272 235172 700284
rect 235224 700272 235230 700324
rect 267642 700272 267648 700324
rect 267700 700312 267706 700324
rect 357434 700312 357440 700324
rect 267700 700284 357440 700312
rect 267700 700272 267706 700284
rect 357434 700272 357440 700284
rect 357492 700272 357498 700324
rect 374638 700272 374644 700324
rect 374696 700312 374702 700324
rect 397454 700312 397460 700324
rect 374696 700284 397460 700312
rect 374696 700272 374702 700284
rect 397454 700272 397460 700284
rect 397512 700272 397518 700324
rect 431218 700272 431224 700324
rect 431276 700312 431282 700324
rect 462314 700312 462320 700324
rect 431276 700284 462320 700312
rect 431276 700272 431282 700284
rect 462314 700272 462320 700284
rect 462372 700272 462378 700324
rect 462958 700272 462964 700324
rect 463016 700312 463022 700324
rect 559650 700312 559656 700324
rect 463016 700284 559656 700312
rect 463016 700272 463022 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 105446 699728 105452 699780
rect 105504 699768 105510 699780
rect 108298 699768 108304 699780
rect 105504 699740 108304 699768
rect 105504 699728 105510 699740
rect 108298 699728 108304 699740
rect 108356 699728 108362 699780
rect 428458 699660 428464 699712
rect 428516 699700 428522 699712
rect 429838 699700 429844 699712
rect 428516 699672 429844 699700
rect 428516 699660 428522 699672
rect 429838 699660 429844 699672
rect 429896 699660 429902 699712
rect 387058 696940 387064 696992
rect 387116 696980 387122 696992
rect 580166 696980 580172 696992
rect 387116 696952 580172 696980
rect 387116 696940 387122 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 171778 683176 171784 683188
rect 3476 683148 171784 683176
rect 3476 683136 3482 683148
rect 171778 683136 171784 683148
rect 171836 683136 171842 683188
rect 371878 670692 371884 670744
rect 371936 670732 371942 670744
rect 580166 670732 580172 670744
rect 371936 670704 580172 670732
rect 371936 670692 371942 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 21358 656928 21364 656940
rect 3568 656900 21364 656928
rect 3568 656888 3574 656900
rect 21358 656888 21364 656900
rect 21416 656888 21422 656940
rect 373258 643084 373264 643136
rect 373316 643124 373322 643136
rect 580166 643124 580172 643136
rect 373316 643096 580172 643124
rect 373316 643084 373322 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4798 632108 4804 632120
rect 2832 632080 4804 632108
rect 2832 632068 2838 632080
rect 4798 632068 4804 632080
rect 4856 632068 4862 632120
rect 367738 630640 367744 630692
rect 367796 630680 367802 630692
rect 579982 630680 579988 630692
rect 367796 630652 579988 630680
rect 367796 630640 367802 630652
rect 579982 630640 579988 630652
rect 580040 630640 580046 630692
rect 363598 616836 363604 616888
rect 363656 616876 363662 616888
rect 580166 616876 580172 616888
rect 363656 616848 580172 616876
rect 363656 616836 363662 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3326 605820 3332 605872
rect 3384 605860 3390 605872
rect 17218 605860 17224 605872
rect 3384 605832 17224 605860
rect 3384 605820 3390 605832
rect 17218 605820 17224 605832
rect 17276 605820 17282 605872
rect 369118 590656 369124 590708
rect 369176 590696 369182 590708
rect 580166 590696 580172 590708
rect 369176 590668 580172 590696
rect 369176 590656 369182 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 10318 579680 10324 579692
rect 3384 579652 10324 579680
rect 3384 579640 3390 579652
rect 10318 579640 10324 579652
rect 10376 579640 10382 579692
rect 359458 576852 359464 576904
rect 359516 576892 359522 576904
rect 580166 576892 580172 576904
rect 359516 576864 580172 576892
rect 359516 576852 359522 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3142 553664 3148 553716
rect 3200 553704 3206 553716
rect 8938 553704 8944 553716
rect 3200 553676 8944 553704
rect 3200 553664 3206 553676
rect 8938 553664 8944 553676
rect 8996 553664 9002 553716
rect 3326 527144 3332 527196
rect 3384 527184 3390 527196
rect 14458 527184 14464 527196
rect 3384 527156 14464 527184
rect 3384 527144 3390 527156
rect 14458 527144 14464 527156
rect 14516 527144 14522 527196
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 18598 514808 18604 514820
rect 3384 514780 18604 514808
rect 3384 514768 3390 514780
rect 18598 514768 18604 514780
rect 18656 514768 18662 514820
rect 2866 500964 2872 501016
rect 2924 501004 2930 501016
rect 13078 501004 13084 501016
rect 2924 500976 13084 501004
rect 2924 500964 2930 500976
rect 13078 500964 13084 500976
rect 13136 500964 13142 501016
rect 360838 563048 360844 563100
rect 360896 563088 360902 563100
rect 580166 563088 580172 563100
rect 360896 563060 580172 563088
rect 360896 563048 360902 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 496078 536800 496084 536852
rect 496136 536840 496142 536852
rect 579890 536840 579896 536852
rect 496136 536812 579896 536840
rect 496136 536800 496142 536812
rect 579890 536800 579896 536812
rect 579948 536800 579954 536852
rect 480898 484372 480904 484424
rect 480956 484412 480962 484424
rect 580166 484412 580172 484424
rect 480956 484384 580172 484412
rect 480956 484372 480962 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 217318 478864 217324 478916
rect 217376 478904 217382 478916
rect 220078 478904 220084 478916
rect 217376 478876 220084 478904
rect 217376 478864 217382 478876
rect 220078 478864 220084 478876
rect 220136 478864 220142 478916
rect 309134 478252 309140 478304
rect 309192 478292 309198 478304
rect 357710 478292 357716 478304
rect 309192 478264 357716 478292
rect 309192 478252 309198 478264
rect 357710 478252 357716 478264
rect 357768 478252 357774 478304
rect 218054 478184 218060 478236
rect 218112 478224 218118 478236
rect 313366 478224 313372 478236
rect 218112 478196 313372 478224
rect 218112 478184 218118 478196
rect 313366 478184 313372 478196
rect 313424 478184 313430 478236
rect 21358 478116 21364 478168
rect 21416 478156 21422 478168
rect 346486 478156 346492 478168
rect 21416 478128 346492 478156
rect 21416 478116 21422 478128
rect 346486 478116 346492 478128
rect 346544 478116 346550 478168
rect 217502 476756 217508 476808
rect 217560 476796 217566 476808
rect 233326 476796 233332 476808
rect 217560 476768 233332 476796
rect 217560 476756 217566 476768
rect 233326 476756 233332 476768
rect 233384 476756 233390 476808
rect 255406 476756 255412 476808
rect 255464 476796 255470 476808
rect 264974 476796 264980 476808
rect 255464 476768 264980 476796
rect 255464 476756 255470 476768
rect 264974 476756 264980 476768
rect 265032 476756 265038 476808
rect 251174 476688 251180 476740
rect 251232 476728 251238 476740
rect 260834 476728 260840 476740
rect 251232 476700 260840 476728
rect 251232 476688 251238 476700
rect 260834 476688 260840 476700
rect 260892 476688 260898 476740
rect 277578 476688 277584 476740
rect 277636 476728 277642 476740
rect 302234 476728 302240 476740
rect 277636 476700 302240 476728
rect 277636 476688 277642 476700
rect 302234 476688 302240 476700
rect 302292 476688 302298 476740
rect 255222 476620 255228 476672
rect 255280 476660 255286 476672
rect 259454 476660 259460 476672
rect 255280 476632 259460 476660
rect 255280 476620 255286 476632
rect 259454 476620 259460 476632
rect 259512 476620 259518 476672
rect 278774 476620 278780 476672
rect 278832 476660 278838 476672
rect 304994 476660 305000 476672
rect 278832 476632 305000 476660
rect 278832 476620 278838 476632
rect 304994 476620 305000 476632
rect 305052 476620 305058 476672
rect 238754 476552 238760 476604
rect 238812 476592 238818 476604
rect 244274 476592 244280 476604
rect 238812 476564 244280 476592
rect 238812 476552 238818 476564
rect 244274 476552 244280 476564
rect 244332 476552 244338 476604
rect 252554 476592 252560 476604
rect 244384 476564 252560 476592
rect 235994 476484 236000 476536
rect 236052 476524 236058 476536
rect 242894 476524 242900 476536
rect 236052 476496 242900 476524
rect 236052 476484 236058 476496
rect 242894 476484 242900 476496
rect 242952 476484 242958 476536
rect 242986 476484 242992 476536
rect 243044 476524 243050 476536
rect 244384 476524 244412 476564
rect 252554 476552 252560 476564
rect 252612 476552 252618 476604
rect 252646 476552 252652 476604
rect 252704 476592 252710 476604
rect 263594 476592 263600 476604
rect 252704 476564 263600 476592
rect 252704 476552 252710 476564
rect 263594 476552 263600 476564
rect 263652 476552 263658 476604
rect 282914 476552 282920 476604
rect 282972 476592 282978 476604
rect 310514 476592 310520 476604
rect 282972 476564 310520 476592
rect 282972 476552 282978 476564
rect 310514 476552 310520 476564
rect 310572 476552 310578 476604
rect 243044 476496 244412 476524
rect 243044 476484 243050 476496
rect 248414 476484 248420 476536
rect 248472 476524 248478 476536
rect 258258 476524 258264 476536
rect 248472 476496 258264 476524
rect 248472 476484 248478 476496
rect 258258 476484 258264 476496
rect 258316 476484 258322 476536
rect 262306 476484 262312 476536
rect 262364 476524 262370 476536
rect 276014 476524 276020 476536
rect 262364 476496 276020 476524
rect 262364 476484 262370 476496
rect 276014 476484 276020 476496
rect 276072 476484 276078 476536
rect 280154 476484 280160 476536
rect 280212 476524 280218 476536
rect 307754 476524 307760 476536
rect 280212 476496 307760 476524
rect 280212 476484 280218 476496
rect 307754 476484 307760 476496
rect 307812 476484 307818 476536
rect 236086 476416 236092 476468
rect 236144 476456 236150 476468
rect 247034 476456 247040 476468
rect 236144 476428 247040 476456
rect 236144 476416 236150 476428
rect 247034 476416 247040 476428
rect 247092 476416 247098 476468
rect 256786 476416 256792 476468
rect 256844 476456 256850 476468
rect 267918 476456 267924 476468
rect 256844 476428 267924 476456
rect 256844 476416 256850 476428
rect 267918 476416 267924 476428
rect 267976 476416 267982 476468
rect 285674 476416 285680 476468
rect 285732 476456 285738 476468
rect 314654 476456 314660 476468
rect 285732 476428 314660 476456
rect 285732 476416 285738 476428
rect 314654 476416 314660 476428
rect 314712 476416 314718 476468
rect 245746 476348 245752 476400
rect 245804 476388 245810 476400
rect 255314 476388 255320 476400
rect 245804 476360 255320 476388
rect 245804 476348 245810 476360
rect 255314 476348 255320 476360
rect 255372 476348 255378 476400
rect 258074 476348 258080 476400
rect 258132 476388 258138 476400
rect 260098 476388 260104 476400
rect 258132 476360 260104 476388
rect 258132 476348 258138 476360
rect 260098 476348 260104 476360
rect 260156 476348 260162 476400
rect 260926 476348 260932 476400
rect 260984 476388 260990 476400
rect 273254 476388 273260 476400
rect 260984 476360 273260 476388
rect 260984 476348 260990 476360
rect 273254 476348 273260 476360
rect 273312 476348 273318 476400
rect 284294 476348 284300 476400
rect 284352 476388 284358 476400
rect 313274 476388 313280 476400
rect 284352 476360 313280 476388
rect 284352 476348 284358 476360
rect 313274 476348 313280 476360
rect 313332 476348 313338 476400
rect 237282 476280 237288 476332
rect 237340 476320 237346 476332
rect 238846 476320 238852 476332
rect 237340 476292 238852 476320
rect 237340 476280 237346 476292
rect 238846 476280 238852 476292
rect 238904 476280 238910 476332
rect 240134 476280 240140 476332
rect 240192 476320 240198 476332
rect 240192 476292 248414 476320
rect 240192 476280 240198 476292
rect 241514 476212 241520 476264
rect 241572 476252 241578 476264
rect 244274 476252 244280 476264
rect 241572 476224 244280 476252
rect 241572 476212 241578 476224
rect 244274 476212 244280 476224
rect 244332 476212 244338 476264
rect 248386 476252 248414 476292
rect 258166 476280 258172 476332
rect 258224 476320 258230 476332
rect 258224 476292 267734 476320
rect 258224 476280 258230 476292
rect 249886 476252 249892 476264
rect 248386 476224 249892 476252
rect 249886 476212 249892 476224
rect 249944 476212 249950 476264
rect 263686 476212 263692 476264
rect 263744 476252 263750 476264
rect 267706 476252 267734 476292
rect 287054 476280 287060 476332
rect 287112 476320 287118 476332
rect 317414 476320 317420 476332
rect 287112 476292 317420 476320
rect 287112 476280 287118 476292
rect 317414 476280 317420 476292
rect 317472 476280 317478 476332
rect 270494 476252 270500 476264
rect 263744 476224 264376 476252
rect 267706 476224 270500 476252
rect 263744 476212 263750 476224
rect 242802 476144 242808 476196
rect 242860 476184 242866 476196
rect 244918 476184 244924 476196
rect 242860 476156 244924 476184
rect 242860 476144 242866 476156
rect 244918 476144 244924 476156
rect 244976 476144 244982 476196
rect 262122 476144 262128 476196
rect 262180 476184 262186 476196
rect 264238 476184 264244 476196
rect 262180 476156 264244 476184
rect 262180 476144 262186 476156
rect 264238 476144 264244 476156
rect 264296 476144 264302 476196
rect 264348 476184 264376 476224
rect 270494 476212 270500 476224
rect 270552 476212 270558 476264
rect 288434 476212 288440 476264
rect 288492 476252 288498 476264
rect 320174 476252 320180 476264
rect 288492 476224 320180 476252
rect 288492 476212 288498 476224
rect 320174 476212 320180 476224
rect 320232 476212 320238 476264
rect 264348 476156 267734 476184
rect 234614 476076 234620 476128
rect 234672 476116 234678 476128
rect 235902 476116 235908 476128
rect 234672 476088 235908 476116
rect 234672 476076 234678 476088
rect 235902 476076 235908 476088
rect 235960 476076 235966 476128
rect 241422 476076 241428 476128
rect 241480 476116 241486 476128
rect 242986 476116 242992 476128
rect 241480 476088 242992 476116
rect 241480 476076 241486 476088
rect 242986 476076 242992 476088
rect 243044 476076 243050 476128
rect 244274 476076 244280 476128
rect 244332 476116 244338 476128
rect 245654 476116 245660 476128
rect 244332 476088 245660 476116
rect 244332 476076 244338 476088
rect 245654 476076 245660 476088
rect 245712 476076 245718 476128
rect 252462 476076 252468 476128
rect 252520 476116 252526 476128
rect 253934 476116 253940 476128
rect 252520 476088 253940 476116
rect 252520 476076 252526 476088
rect 253934 476076 253940 476088
rect 253992 476076 253998 476128
rect 260742 476076 260748 476128
rect 260800 476116 260806 476128
rect 262858 476116 262864 476128
rect 260800 476088 262864 476116
rect 260800 476076 260806 476088
rect 262858 476076 262864 476088
rect 262916 476076 262922 476128
rect 263502 476076 263508 476128
rect 263560 476116 263566 476128
rect 265618 476116 265624 476128
rect 263560 476088 265624 476116
rect 263560 476076 263566 476088
rect 265618 476076 265624 476088
rect 265676 476076 265682 476128
rect 267706 476116 267734 476156
rect 289814 476144 289820 476196
rect 289872 476184 289878 476196
rect 322934 476184 322940 476196
rect 289872 476156 322940 476184
rect 289872 476144 289878 476156
rect 322934 476144 322940 476156
rect 322992 476144 322998 476196
rect 277854 476116 277860 476128
rect 267706 476088 277860 476116
rect 277854 476076 277860 476088
rect 277912 476076 277918 476128
rect 291194 476076 291200 476128
rect 291252 476116 291258 476128
rect 325786 476116 325792 476128
rect 291252 476088 325792 476116
rect 291252 476076 291258 476088
rect 325786 476076 325792 476088
rect 325844 476076 325850 476128
rect 219066 475328 219072 475380
rect 219124 475368 219130 475380
rect 241606 475368 241612 475380
rect 219124 475340 241612 475368
rect 219124 475328 219130 475340
rect 241606 475328 241612 475340
rect 241664 475328 241670 475380
rect 302234 475328 302240 475380
rect 302292 475368 302298 475380
rect 542354 475368 542360 475380
rect 302292 475340 542360 475368
rect 302292 475328 302298 475340
rect 542354 475328 542360 475340
rect 542412 475328 542418 475380
rect 3326 474716 3332 474768
rect 3384 474756 3390 474768
rect 329834 474756 329840 474768
rect 3384 474728 329840 474756
rect 3384 474716 3390 474728
rect 329834 474716 329840 474728
rect 329892 474716 329898 474768
rect 219158 474036 219164 474088
rect 219216 474076 219222 474088
rect 247126 474076 247132 474088
rect 219216 474048 247132 474076
rect 219216 474036 219222 474048
rect 247126 474036 247132 474048
rect 247184 474036 247190 474088
rect 6914 473968 6920 474020
rect 6972 474008 6978 474020
rect 345106 474008 345112 474020
rect 6972 473980 345112 474008
rect 6972 473968 6978 473980
rect 345106 473968 345112 473980
rect 345164 473968 345170 474020
rect 217686 472676 217692 472728
rect 217744 472716 217750 472728
rect 251266 472716 251272 472728
rect 217744 472688 251272 472716
rect 217744 472676 217750 472688
rect 251266 472676 251272 472688
rect 251324 472676 251330 472728
rect 332594 472676 332600 472728
rect 332652 472716 332658 472728
rect 374638 472716 374644 472728
rect 332652 472688 374644 472716
rect 332652 472676 332658 472688
rect 374638 472676 374644 472688
rect 374696 472676 374702 472728
rect 17218 472608 17224 472660
rect 17276 472648 17282 472660
rect 347774 472648 347780 472660
rect 17276 472620 347780 472648
rect 17276 472608 17282 472620
rect 347774 472608 347780 472620
rect 347832 472608 347838 472660
rect 217778 471316 217784 471368
rect 217836 471356 217842 471368
rect 254026 471356 254032 471368
rect 217836 471328 254032 471356
rect 217836 471316 217842 471328
rect 254026 471316 254032 471328
rect 254084 471316 254090 471368
rect 299474 471316 299480 471368
rect 299532 471356 299538 471368
rect 580258 471356 580264 471368
rect 299532 471328 580264 471356
rect 299532 471316 299538 471328
rect 580258 471316 580264 471328
rect 580316 471316 580322 471368
rect 14458 471248 14464 471300
rect 14516 471288 14522 471300
rect 327074 471288 327080 471300
rect 14516 471260 327080 471288
rect 14516 471248 14522 471260
rect 327074 471248 327080 471260
rect 327132 471248 327138 471300
rect 267826 469888 267832 469940
rect 267884 469928 267890 469940
rect 285766 469928 285772 469940
rect 267884 469900 285772 469928
rect 267884 469888 267890 469900
rect 285766 469888 285772 469900
rect 285824 469888 285830 469940
rect 298094 469888 298100 469940
rect 298152 469928 298158 469940
rect 367738 469928 367744 469940
rect 298152 469900 367744 469928
rect 298152 469888 298158 469900
rect 367738 469888 367744 469900
rect 367796 469888 367802 469940
rect 10318 469820 10324 469872
rect 10376 469860 10382 469872
rect 324314 469860 324320 469872
rect 10376 469832 324320 469860
rect 10376 469820 10382 469832
rect 324314 469820 324320 469832
rect 324372 469820 324378 469872
rect 269206 468528 269212 468580
rect 269264 468568 269270 468580
rect 287146 468568 287152 468580
rect 269264 468540 287152 468568
rect 269264 468528 269270 468540
rect 287146 468528 287152 468540
rect 287204 468528 287210 468580
rect 108298 468460 108304 468512
rect 108356 468500 108362 468512
rect 316034 468500 316040 468512
rect 108356 468472 316040 468500
rect 108356 468460 108362 468472
rect 316034 468460 316040 468472
rect 316092 468460 316098 468512
rect 318794 468460 318800 468512
rect 318852 468500 318858 468512
rect 496078 468500 496084 468512
rect 318852 468472 496084 468500
rect 318852 468460 318858 468472
rect 496078 468460 496084 468472
rect 496136 468460 496142 468512
rect 295334 467168 295340 467220
rect 295392 467208 295398 467220
rect 359458 467208 359464 467220
rect 295392 467180 359464 467208
rect 295392 467168 295398 467180
rect 359458 467168 359464 467180
rect 359516 467168 359522 467220
rect 171778 467100 171784 467152
rect 171836 467140 171842 467152
rect 320174 467140 320180 467152
rect 171836 467112 320180 467140
rect 171836 467100 171842 467112
rect 320174 467100 320180 467112
rect 320232 467100 320238 467152
rect 4798 465672 4804 465724
rect 4856 465712 4862 465724
rect 322934 465712 322940 465724
rect 4856 465684 322940 465712
rect 4856 465672 4862 465684
rect 322934 465672 322940 465684
rect 322992 465672 322998 465724
rect 325694 465672 325700 465724
rect 325752 465712 325758 465724
rect 387058 465712 387064 465724
rect 325752 465684 387064 465712
rect 325752 465672 325758 465684
rect 387058 465672 387064 465684
rect 387116 465672 387122 465724
rect 169754 464312 169760 464364
rect 169812 464352 169818 464364
rect 313366 464352 313372 464364
rect 169812 464324 313372 464352
rect 169812 464312 169818 464324
rect 313366 464312 313372 464324
rect 313424 464312 313430 464364
rect 323026 464312 323032 464364
rect 323084 464352 323090 464364
rect 373258 464352 373264 464364
rect 323084 464324 373264 464352
rect 323084 464312 323090 464324
rect 373258 464312 373264 464324
rect 373316 464312 373322 464364
rect 329926 462952 329932 463004
rect 329984 462992 329990 463004
rect 431218 462992 431224 463004
rect 329984 462964 431224 462992
rect 329984 462952 329990 462964
rect 431218 462952 431224 462964
rect 431276 462952 431282 463004
rect 3326 462340 3332 462392
rect 3384 462380 3390 462392
rect 331306 462380 331312 462392
rect 3384 462352 331312 462380
rect 3384 462340 3390 462352
rect 331306 462340 331312 462352
rect 331364 462340 331370 462392
rect 40034 461592 40040 461644
rect 40092 461632 40098 461644
rect 318886 461632 318892 461644
rect 40092 461604 318892 461632
rect 40092 461592 40098 461604
rect 318886 461592 318892 461604
rect 318944 461592 318950 461644
rect 321554 461592 321560 461644
rect 321612 461632 321618 461644
rect 369118 461632 369124 461644
rect 321612 461604 369124 461632
rect 321612 461592 321618 461604
rect 369118 461592 369124 461604
rect 369176 461592 369182 461644
rect 270770 460232 270776 460284
rect 270828 460272 270834 460284
rect 289906 460272 289912 460284
rect 270828 460244 289912 460272
rect 270828 460232 270834 460244
rect 289906 460232 289912 460244
rect 289964 460232 289970 460284
rect 307754 460232 307760 460284
rect 307812 460272 307818 460284
rect 364334 460272 364340 460284
rect 307812 460244 364340 460272
rect 307812 460232 307818 460244
rect 364334 460232 364340 460244
rect 364392 460232 364398 460284
rect 8938 460164 8944 460216
rect 8996 460204 9002 460216
rect 349154 460204 349160 460216
rect 8996 460176 349160 460204
rect 8996 460164 9002 460176
rect 349154 460164 349160 460176
rect 349212 460164 349218 460216
rect 273162 458872 273168 458924
rect 273220 458912 273226 458924
rect 281810 458912 281816 458924
rect 273220 458884 281816 458912
rect 273220 458872 273226 458884
rect 281810 458872 281816 458884
rect 281868 458872 281874 458924
rect 219250 458804 219256 458856
rect 219308 458844 219314 458856
rect 244366 458844 244372 458856
rect 219308 458816 244372 458844
rect 219308 458804 219314 458816
rect 244366 458804 244372 458816
rect 244424 458804 244430 458856
rect 278682 458804 278688 458856
rect 278740 458844 278746 458856
rect 289170 458844 289176 458856
rect 278740 458816 289176 458844
rect 278740 458804 278746 458816
rect 289170 458804 289176 458816
rect 289228 458804 289234 458856
rect 317414 458804 317420 458856
rect 317472 458844 317478 458856
rect 480898 458844 480904 458856
rect 317472 458816 480904 458844
rect 317472 458804 317478 458816
rect 480898 458804 480904 458816
rect 480956 458804 480962 458856
rect 266446 457512 266452 457564
rect 266504 457552 266510 457564
rect 283006 457552 283012 457564
rect 266504 457524 283012 457552
rect 266504 457512 266510 457524
rect 283006 457512 283012 457524
rect 283064 457512 283070 457564
rect 305362 457512 305368 457564
rect 305420 457552 305426 457564
rect 428458 457552 428464 457564
rect 305420 457524 428464 457552
rect 305420 457512 305426 457524
rect 428458 457512 428464 457524
rect 428516 457512 428522 457564
rect 13078 457444 13084 457496
rect 13136 457484 13142 457496
rect 349522 457484 349528 457496
rect 13136 457456 349528 457484
rect 13136 457444 13142 457456
rect 349522 457444 349528 457456
rect 349580 457444 349586 457496
rect 265066 456084 265072 456136
rect 265124 456124 265130 456136
rect 280246 456124 280252 456136
rect 265124 456096 280252 456124
rect 265124 456084 265130 456096
rect 280246 456084 280252 456096
rect 280304 456084 280310 456136
rect 303154 456084 303160 456136
rect 303212 456124 303218 456136
rect 494054 456124 494060 456136
rect 303212 456096 494060 456124
rect 303212 456084 303218 456096
rect 494054 456084 494060 456096
rect 494112 456084 494118 456136
rect 18598 456016 18604 456068
rect 18656 456056 18662 456068
rect 328914 456056 328920 456068
rect 18656 456028 328920 456056
rect 18656 456016 18662 456028
rect 328914 456016 328920 456028
rect 328972 456016 328978 456068
rect 274450 454792 274456 454844
rect 274508 454832 274514 454844
rect 283282 454832 283288 454844
rect 274508 454804 283288 454832
rect 274508 454792 274514 454804
rect 283282 454792 283288 454804
rect 283340 454792 283346 454844
rect 276014 454724 276020 454776
rect 276072 454764 276078 454776
rect 300854 454764 300860 454776
rect 276072 454736 300860 454764
rect 276072 454724 276078 454736
rect 300854 454724 300860 454736
rect 300912 454724 300918 454776
rect 217870 454656 217876 454708
rect 217928 454696 217934 454708
rect 256050 454696 256056 454708
rect 217928 454668 256056 454696
rect 217928 454656 217934 454668
rect 256050 454656 256056 454668
rect 256108 454656 256114 454708
rect 267550 454656 267556 454708
rect 267608 454696 267614 454708
rect 276106 454696 276112 454708
rect 267608 454668 276112 454696
rect 267608 454656 267614 454668
rect 276106 454656 276112 454668
rect 276164 454656 276170 454708
rect 280062 454656 280068 454708
rect 280120 454696 280126 454708
rect 290642 454696 290648 454708
rect 280120 454668 290648 454696
rect 280120 454656 280126 454668
rect 290642 454656 290648 454668
rect 290700 454656 290706 454708
rect 298738 454656 298744 454708
rect 298796 454696 298802 454708
rect 371878 454696 371884 454708
rect 298796 454668 371884 454696
rect 298796 454656 298802 454668
rect 371878 454656 371884 454668
rect 371936 454656 371942 454708
rect 271782 453432 271788 453484
rect 271840 453472 271846 453484
rect 280338 453472 280344 453484
rect 271840 453444 280344 453472
rect 271840 453432 271846 453444
rect 280338 453432 280344 453444
rect 280396 453432 280402 453484
rect 277302 453364 277308 453416
rect 277360 453404 277366 453416
rect 287698 453404 287704 453416
rect 277360 453376 287704 453404
rect 277360 453364 277366 453376
rect 287698 453364 287704 453376
rect 287756 453364 287762 453416
rect 267642 453296 267648 453348
rect 267700 453336 267706 453348
rect 274634 453336 274640 453348
rect 267700 453308 274640 453336
rect 267700 453296 267706 453308
rect 274634 453296 274640 453308
rect 274692 453296 274698 453348
rect 275186 453296 275192 453348
rect 275244 453336 275250 453348
rect 298186 453336 298192 453348
rect 275244 453308 298192 453336
rect 275244 453296 275250 453308
rect 298186 453296 298192 453308
rect 298244 453296 298250 453348
rect 300946 453296 300952 453348
rect 301004 453336 301010 453348
rect 462958 453336 462964 453348
rect 301004 453308 462964 453336
rect 301004 453296 301010 453308
rect 462958 453296 462964 453308
rect 463016 453296 463022 453348
rect 269022 452004 269028 452056
rect 269080 452044 269086 452056
rect 277486 452044 277492 452056
rect 269080 452016 277492 452044
rect 269080 452004 269086 452016
rect 277486 452004 277492 452016
rect 277544 452004 277550 452056
rect 275922 451936 275928 451988
rect 275980 451976 275986 451988
rect 286226 451976 286232 451988
rect 275980 451948 286232 451976
rect 275980 451936 275986 451948
rect 286226 451936 286232 451948
rect 286284 451936 286290 451988
rect 217594 451868 217600 451920
rect 217652 451908 217658 451920
rect 234706 451908 234712 451920
rect 217652 451880 234712 451908
rect 217652 451868 217658 451880
rect 234706 451868 234712 451880
rect 234764 451868 234770 451920
rect 264882 451868 264888 451920
rect 264940 451908 264946 451920
rect 271874 451908 271880 451920
rect 264940 451880 271880 451908
rect 264940 451868 264946 451880
rect 271874 451868 271880 451880
rect 271932 451868 271938 451920
rect 272242 451868 272248 451920
rect 272300 451908 272306 451920
rect 292574 451908 292580 451920
rect 272300 451880 292580 451908
rect 272300 451868 272306 451880
rect 292574 451868 292580 451880
rect 292632 451868 292638 451920
rect 296714 451868 296720 451920
rect 296772 451908 296778 451920
rect 363598 451908 363604 451920
rect 296772 451880 363604 451908
rect 296772 451868 296778 451880
rect 363598 451868 363604 451880
rect 363656 451868 363662 451920
rect 270402 450644 270408 450696
rect 270460 450684 270466 450696
rect 279234 450684 279240 450696
rect 270460 450656 279240 450684
rect 270460 450644 270466 450656
rect 279234 450644 279240 450656
rect 279292 450644 279298 450696
rect 274082 450576 274088 450628
rect 274140 450616 274146 450628
rect 295426 450616 295432 450628
rect 274140 450588 295432 450616
rect 274140 450576 274146 450588
rect 295426 450576 295432 450588
rect 295484 450576 295490 450628
rect 219342 450508 219348 450560
rect 219400 450548 219406 450560
rect 249794 450548 249800 450560
rect 219400 450520 249800 450548
rect 219400 450508 219406 450520
rect 249794 450508 249800 450520
rect 249852 450508 249858 450560
rect 266262 450508 266268 450560
rect 266320 450548 266326 450560
rect 273346 450548 273352 450560
rect 266320 450520 273352 450548
rect 266320 450508 266326 450520
rect 273346 450508 273352 450520
rect 273404 450508 273410 450560
rect 274542 450508 274548 450560
rect 274600 450548 274606 450560
rect 285122 450548 285128 450560
rect 274600 450520 285128 450548
rect 274600 450508 274606 450520
rect 285122 450508 285128 450520
rect 285180 450508 285186 450560
rect 294690 450508 294696 450560
rect 294748 450548 294754 450560
rect 360838 450548 360844 450560
rect 294748 450520 360844 450548
rect 294748 450508 294754 450520
rect 360838 450508 360844 450520
rect 360896 450508 360902 450560
rect 307202 449624 307208 449676
rect 307260 449664 307266 449676
rect 412634 449664 412640 449676
rect 307260 449636 412640 449664
rect 307260 449624 307266 449636
rect 412634 449624 412640 449636
rect 412692 449624 412698 449676
rect 153194 449556 153200 449608
rect 153252 449596 153258 449608
rect 316034 449596 316040 449608
rect 153252 449568 316040 449596
rect 153252 449556 153258 449568
rect 316034 449556 316040 449568
rect 316092 449556 316098 449608
rect 304994 449488 305000 449540
rect 305052 449528 305058 449540
rect 477494 449528 477500 449540
rect 305052 449500 477500 449528
rect 305052 449488 305058 449500
rect 477494 449488 477500 449500
rect 477552 449488 477558 449540
rect 88334 449420 88340 449472
rect 88392 449460 88398 449472
rect 318242 449460 318248 449472
rect 88392 449432 318248 449460
rect 88392 449420 88398 449432
rect 318242 449420 318248 449432
rect 318300 449420 318306 449472
rect 23474 449352 23480 449404
rect 23532 449392 23538 449404
rect 320450 449392 320456 449404
rect 23532 449364 320456 449392
rect 23532 449352 23538 449364
rect 320450 449352 320456 449364
rect 320508 449352 320514 449404
rect 3418 449284 3424 449336
rect 3476 449324 3482 449336
rect 322658 449324 322664 449336
rect 3476 449296 322664 449324
rect 3476 449284 3482 449296
rect 322658 449284 322664 449296
rect 322716 449284 322722 449336
rect 3510 449216 3516 449268
rect 3568 449256 3574 449268
rect 324866 449256 324872 449268
rect 3568 449228 324872 449256
rect 3568 449216 3574 449228
rect 324866 449216 324872 449228
rect 324924 449216 324930 449268
rect 3602 449148 3608 449200
rect 3660 449188 3666 449200
rect 327074 449188 327080 449200
rect 3660 449160 327080 449188
rect 3660 449148 3666 449160
rect 327074 449148 327080 449160
rect 327132 449148 327138 449200
rect 201494 448060 201500 448112
rect 201552 448100 201558 448112
rect 339586 448100 339592 448112
rect 201552 448072 339592 448100
rect 201552 448060 201558 448072
rect 339586 448060 339592 448072
rect 339644 448060 339650 448112
rect 328546 447992 328552 448044
rect 328604 448032 328610 448044
rect 527174 448032 527180 448044
rect 328604 448004 527180 448032
rect 328604 447992 328610 448004
rect 527174 447992 527180 448004
rect 527232 447992 527238 448044
rect 136634 447924 136640 447976
rect 136692 447964 136698 447976
rect 341794 447964 341800 447976
rect 136692 447936 341800 447964
rect 136692 447924 136698 447936
rect 341794 447924 341800 447936
rect 341852 447924 341858 447976
rect 71774 447856 71780 447908
rect 71832 447896 71838 447908
rect 344002 447896 344008 447908
rect 71832 447868 344008 447896
rect 71832 447856 71838 447868
rect 344002 447856 344008 447868
rect 344060 447856 344066 447908
rect 2866 447788 2872 447840
rect 2924 447828 2930 447840
rect 350626 447828 350632 447840
rect 2924 447800 350632 447828
rect 2924 447788 2930 447800
rect 350626 447788 350632 447800
rect 350684 447788 350690 447840
rect 254578 447040 254584 447092
rect 254636 447080 254642 447092
rect 258626 447080 258632 447092
rect 254636 447052 258632 447080
rect 254636 447040 254642 447052
rect 258626 447040 258632 447052
rect 258684 447040 258690 447092
rect 262858 447040 262864 447092
rect 262916 447080 262922 447092
rect 267458 447080 267464 447092
rect 262916 447052 267464 447080
rect 262916 447040 262922 447052
rect 267458 447040 267464 447052
rect 267516 447040 267522 447092
rect 270402 447080 270408 447092
rect 267706 447052 270408 447080
rect 234614 446972 234620 447024
rect 234672 447012 234678 447024
rect 235534 447012 235540 447024
rect 234672 446984 235540 447012
rect 234672 446972 234678 446984
rect 235534 446972 235540 446984
rect 235592 446972 235598 447024
rect 238754 446972 238760 447024
rect 238812 447012 238818 447024
rect 239214 447012 239220 447024
rect 238812 446984 239220 447012
rect 238812 446972 238818 446984
rect 239214 446972 239220 446984
rect 239272 446972 239278 447024
rect 241514 446972 241520 447024
rect 241572 447012 241578 447024
rect 242158 447012 242164 447024
rect 241572 446984 242164 447012
rect 241572 446972 241578 446984
rect 242158 446972 242164 446984
rect 242216 446972 242222 447024
rect 244274 446972 244280 447024
rect 244332 447012 244338 447024
rect 245102 447012 245108 447024
rect 244332 446984 245108 447012
rect 244332 446972 244338 446984
rect 245102 446972 245108 446984
rect 245160 446972 245166 447024
rect 251818 446972 251824 447024
rect 251876 447012 251882 447024
rect 252738 447012 252744 447024
rect 251876 446984 252744 447012
rect 251876 446972 251882 446984
rect 252738 446972 252744 446984
rect 252796 446972 252802 447024
rect 253934 446972 253940 447024
rect 253992 447012 253998 447024
rect 254670 447012 254676 447024
rect 253992 446984 254676 447012
rect 253992 446972 253998 446984
rect 254670 446972 254676 446984
rect 254728 446972 254734 447024
rect 261478 446972 261484 447024
rect 261536 447012 261542 447024
rect 265986 447012 265992 447024
rect 261536 446984 265992 447012
rect 261536 446972 261542 446984
rect 265986 446972 265992 446984
rect 266044 446972 266050 447024
rect 267706 447012 267734 447052
rect 270402 447040 270408 447052
rect 270460 447040 270466 447092
rect 266096 446984 267734 447012
rect 260098 446904 260104 446956
rect 260156 446944 260162 446956
rect 264514 446944 264520 446956
rect 260156 446916 264520 446944
rect 260156 446904 260162 446916
rect 264514 446904 264520 446916
rect 264572 446904 264578 446956
rect 265618 446904 265624 446956
rect 265676 446944 265682 446956
rect 266096 446944 266124 446984
rect 276014 446972 276020 447024
rect 276072 447012 276078 447024
rect 276750 447012 276756 447024
rect 276072 446984 276756 447012
rect 276072 446972 276078 446984
rect 276750 446972 276756 446984
rect 276808 446972 276814 447024
rect 280154 446972 280160 447024
rect 280212 447012 280218 447024
rect 281166 447012 281172 447024
rect 280212 446984 281172 447012
rect 280212 446972 280218 446984
rect 281166 446972 281172 446984
rect 281224 446972 281230 447024
rect 268930 446944 268936 446956
rect 265676 446916 266124 446944
rect 267706 446916 268936 446944
rect 265676 446904 265682 446916
rect 264238 446836 264244 446888
rect 264296 446876 264302 446888
rect 267706 446876 267734 446916
rect 268930 446904 268936 446916
rect 268988 446904 268994 446956
rect 264296 446848 267734 446876
rect 264296 446836 264302 446848
rect 217962 446700 217968 446752
rect 218020 446740 218026 446752
rect 312354 446740 312360 446752
rect 218020 446712 312360 446740
rect 218020 446700 218026 446712
rect 312354 446700 312360 446712
rect 312412 446700 312418 446752
rect 335170 446632 335176 446684
rect 335228 446672 335234 446684
rect 358814 446672 358820 446684
rect 335228 446644 358820 446672
rect 335228 446632 335234 446644
rect 358814 446632 358820 446644
rect 358872 446632 358878 446684
rect 302050 446564 302056 446616
rect 302108 446604 302114 446616
rect 333974 446604 333980 446616
rect 302108 446576 333980 446604
rect 302108 446564 302114 446576
rect 333974 446564 333980 446576
rect 334032 446564 334038 446616
rect 337378 446564 337384 446616
rect 337436 446604 337442 446616
rect 357434 446604 357440 446616
rect 337436 446576 357440 446604
rect 337436 446564 337442 446576
rect 357434 446564 357440 446576
rect 357492 446564 357498 446616
rect 253198 446496 253204 446548
rect 253256 446536 253262 446548
rect 257154 446536 257160 446548
rect 253256 446508 257160 446536
rect 253256 446496 253262 446508
rect 257154 446496 257160 446508
rect 257212 446496 257218 446548
rect 257982 446496 257988 446548
rect 258040 446536 258046 446548
rect 263042 446536 263048 446548
rect 258040 446508 263048 446536
rect 258040 446496 258046 446508
rect 263042 446496 263048 446508
rect 263100 446496 263106 446548
rect 311618 446496 311624 446548
rect 311676 446536 311682 446548
rect 357526 446536 357532 446548
rect 311676 446508 357532 446536
rect 311676 446496 311682 446508
rect 357526 446496 357532 446508
rect 357584 446496 357590 446548
rect 220078 446428 220084 446480
rect 220136 446468 220142 446480
rect 234338 446468 234344 446480
rect 220136 446440 234344 446468
rect 220136 446428 220142 446440
rect 234338 446428 234344 446440
rect 234396 446428 234402 446480
rect 256602 446428 256608 446480
rect 256660 446468 256666 446480
rect 261570 446468 261576 446480
rect 256660 446440 261576 446468
rect 256660 446428 256666 446440
rect 261570 446428 261576 446440
rect 261628 446428 261634 446480
rect 310146 446428 310152 446480
rect 310204 446468 310210 446480
rect 357618 446468 357624 446480
rect 310204 446440 357624 446468
rect 310204 446428 310210 446440
rect 357618 446428 357624 446440
rect 357676 446428 357682 446480
rect 310882 446360 310888 446412
rect 310940 446400 310946 446412
rect 362218 446400 362224 446412
rect 310940 446372 362224 446400
rect 310940 446360 310946 446372
rect 362218 446360 362224 446372
rect 362276 446360 362282 446412
rect 306466 446292 306472 446344
rect 306524 446332 306530 446344
rect 363598 446332 363604 446344
rect 306524 446304 363604 446332
rect 306524 446292 306530 446304
rect 363598 446292 363604 446304
rect 363656 446292 363662 446344
rect 244918 446224 244924 446276
rect 244976 446264 244982 446276
rect 246850 446264 246856 446276
rect 244976 446236 246856 446264
rect 244976 446224 244982 446236
rect 246850 446224 246856 446236
rect 246908 446224 246914 446276
rect 304258 446224 304264 446276
rect 304316 446264 304322 446276
rect 360838 446264 360844 446276
rect 304316 446236 360844 446264
rect 304316 446224 304322 446236
rect 360838 446224 360844 446236
rect 360896 446224 360902 446276
rect 293218 446156 293224 446208
rect 293276 446196 293282 446208
rect 359458 446196 359464 446208
rect 293276 446168 359464 446196
rect 293276 446156 293282 446168
rect 359458 446156 359464 446168
rect 359516 446156 359522 446208
rect 292482 446088 292488 446140
rect 292540 446128 292546 446140
rect 373258 446128 373264 446140
rect 292540 446100 373264 446128
rect 292540 446088 292546 446100
rect 373258 446088 373264 446100
rect 373316 446088 373322 446140
rect 251082 446020 251088 446072
rect 251140 446060 251146 446072
rect 342530 446060 342536 446072
rect 251140 446032 342536 446060
rect 251140 446020 251146 446032
rect 342530 446020 342536 446032
rect 342588 446020 342594 446072
rect 230934 445952 230940 446004
rect 230992 445992 230998 446004
rect 335906 445992 335912 446004
rect 230992 445964 335912 445992
rect 230992 445952 230998 445964
rect 335906 445952 335912 445964
rect 335964 445952 335970 446004
rect 229738 445884 229744 445936
rect 229796 445924 229802 445936
rect 344738 445924 344744 445936
rect 229796 445896 344744 445924
rect 229796 445884 229802 445896
rect 344738 445884 344744 445896
rect 344796 445884 344802 445936
rect 293954 445816 293960 445868
rect 294012 445856 294018 445868
rect 454678 445856 454684 445868
rect 294012 445828 454684 445856
rect 294012 445816 294018 445828
rect 454678 445816 454684 445828
rect 454736 445816 454742 445868
rect 10318 445748 10324 445800
rect 10376 445788 10382 445800
rect 346946 445788 346952 445800
rect 10376 445760 346952 445788
rect 10376 445748 10382 445760
rect 346946 445748 346952 445760
rect 347004 445748 347010 445800
rect 228450 445136 228456 445188
rect 228508 445176 228514 445188
rect 336642 445176 336648 445188
rect 228508 445148 336648 445176
rect 228508 445136 228514 445148
rect 336642 445136 336648 445148
rect 336700 445136 336706 445188
rect 229922 445068 229928 445120
rect 229980 445108 229986 445120
rect 334434 445108 334440 445120
rect 229980 445080 334440 445108
rect 229980 445068 229986 445080
rect 334434 445068 334440 445080
rect 334492 445068 334498 445120
rect 318794 445000 318800 445052
rect 318852 445040 318858 445052
rect 319438 445040 319444 445052
rect 318852 445012 319444 445040
rect 318852 445000 318858 445012
rect 319438 445000 319444 445012
rect 319496 445000 319502 445052
rect 333974 445000 333980 445052
rect 334032 445040 334038 445052
rect 580258 445040 580264 445052
rect 334032 445012 580264 445040
rect 334032 445000 334038 445012
rect 580258 445000 580264 445012
rect 580316 445000 580322 445052
rect 225598 444932 225604 444984
rect 225656 444972 225662 444984
rect 338850 444972 338856 444984
rect 225656 444944 338856 444972
rect 225656 444932 225662 444944
rect 338850 444932 338856 444944
rect 338908 444932 338914 444984
rect 230014 444864 230020 444916
rect 230072 444904 230078 444916
rect 351362 444904 351368 444916
rect 230072 444876 351368 444904
rect 230072 444864 230078 444876
rect 351362 444864 351368 444876
rect 351420 444864 351426 444916
rect 224218 444796 224224 444848
rect 224276 444836 224282 444848
rect 352834 444836 352840 444848
rect 224276 444808 352840 444836
rect 224276 444796 224282 444808
rect 352834 444796 352840 444808
rect 352892 444796 352898 444848
rect 295426 444728 295432 444780
rect 295484 444768 295490 444780
rect 494698 444768 494704 444780
rect 295484 444740 494704 444768
rect 295484 444728 295490 444740
rect 494698 444728 494704 444740
rect 494756 444728 494762 444780
rect 95970 444660 95976 444712
rect 96028 444700 96034 444712
rect 341058 444700 341064 444712
rect 96028 444672 341064 444700
rect 96028 444660 96034 444672
rect 341058 444660 341064 444672
rect 341116 444660 341122 444712
rect 93118 444592 93124 444644
rect 93176 444632 93182 444644
rect 343266 444632 343272 444644
rect 93176 444604 343272 444632
rect 93176 444592 93182 444604
rect 343266 444592 343272 444604
rect 343324 444592 343330 444644
rect 86218 444524 86224 444576
rect 86276 444564 86282 444576
rect 345474 444564 345480 444576
rect 86276 444536 345480 444564
rect 86276 444524 86282 444536
rect 345474 444524 345480 444536
rect 345532 444524 345538 444576
rect 84838 444456 84844 444508
rect 84896 444496 84902 444508
rect 355042 444496 355048 444508
rect 84896 444468 355048 444496
rect 84896 444456 84902 444468
rect 355042 444456 355048 444468
rect 355100 444456 355106 444508
rect 7558 444388 7564 444440
rect 7616 444428 7622 444440
rect 332226 444428 332232 444440
rect 7616 444400 332232 444428
rect 7616 444388 7622 444400
rect 332226 444388 332232 444400
rect 332284 444388 332290 444440
rect 315298 443708 315304 443760
rect 315356 443748 315362 443760
rect 360930 443748 360936 443760
rect 315356 443720 360936 443748
rect 315356 443708 315362 443720
rect 360930 443708 360936 443720
rect 360988 443708 360994 443760
rect 3510 443640 3516 443692
rect 3568 443680 3574 443692
rect 251082 443680 251088 443692
rect 3568 443652 251088 443680
rect 3568 443640 3574 443652
rect 251082 443640 251088 443652
rect 251140 443640 251146 443692
rect 313090 443640 313096 443692
rect 313148 443680 313154 443692
rect 367738 443680 367744 443692
rect 313148 443652 367744 443680
rect 313148 443640 313154 443652
rect 367738 443640 367744 443652
rect 367796 443640 367802 443692
rect 308674 443572 308680 443624
rect 308732 443612 308738 443624
rect 364978 443612 364984 443624
rect 308732 443584 364984 443612
rect 308732 443572 308738 443584
rect 364978 443572 364984 443584
rect 365036 443572 365042 443624
rect 228542 443504 228548 443556
rect 228600 443544 228606 443556
rect 333698 443544 333704 443556
rect 228600 443516 333704 443544
rect 228600 443504 228606 443516
rect 333698 443504 333704 443516
rect 333756 443504 333762 443556
rect 228358 443436 228364 443488
rect 228416 443476 228422 443488
rect 338206 443476 338212 443488
rect 228416 443448 338212 443476
rect 228416 443436 228422 443448
rect 338206 443436 338212 443448
rect 338264 443436 338270 443488
rect 229830 443368 229836 443420
rect 229888 443408 229894 443420
rect 351914 443408 351920 443420
rect 229888 443380 351920 443408
rect 229888 443368 229894 443380
rect 351914 443368 351920 443380
rect 351972 443368 351978 443420
rect 300118 443300 300124 443352
rect 300176 443340 300182 443352
rect 442258 443340 442264 443352
rect 300176 443312 442264 443340
rect 300176 443300 300182 443312
rect 442258 443300 442264 443312
rect 442316 443300 442322 443352
rect 157978 443232 157984 443284
rect 158036 443272 158042 443284
rect 340046 443272 340052 443284
rect 158036 443244 340052 443272
rect 158036 443232 158042 443244
rect 340046 443232 340052 443244
rect 340104 443232 340110 443284
rect 97258 443164 97264 443216
rect 97316 443204 97322 443216
rect 353294 443204 353300 443216
rect 97316 443176 353300 443204
rect 97316 443164 97322 443176
rect 353294 443164 353300 443176
rect 353352 443164 353358 443216
rect 95878 443096 95884 443148
rect 95936 443136 95942 443148
rect 355502 443136 355508 443148
rect 95936 443108 355508 443136
rect 95936 443096 95942 443108
rect 355502 443096 355508 443108
rect 355560 443096 355566 443148
rect 94498 443028 94504 443080
rect 94556 443068 94562 443080
rect 354030 443068 354036 443080
rect 94556 443040 354036 443068
rect 94556 443028 94562 443040
rect 354030 443028 354036 443040
rect 354088 443028 354094 443080
rect 14458 442960 14464 443012
rect 14516 443000 14522 443012
rect 356974 443000 356980 443012
rect 14516 442972 356980 443000
rect 14516 442960 14522 442972
rect 356974 442960 356980 442972
rect 357032 442960 357038 443012
rect 3418 442212 3424 442264
rect 3476 442252 3482 442264
rect 230842 442252 230848 442264
rect 3476 442224 230848 442252
rect 3476 442212 3482 442224
rect 230842 442212 230848 442224
rect 230900 442212 230906 442264
rect 359458 442212 359464 442264
rect 359516 442252 359522 442264
rect 580994 442252 581000 442264
rect 359516 442224 581000 442252
rect 359516 442212 359522 442224
rect 580994 442212 581000 442224
rect 581052 442212 581058 442264
rect 3602 440852 3608 440904
rect 3660 440892 3666 440904
rect 230934 440892 230940 440904
rect 3660 440864 230940 440892
rect 3660 440852 3666 440864
rect 230934 440852 230940 440864
rect 230992 440852 230998 440904
rect 454678 438132 454684 438184
rect 454736 438172 454742 438184
rect 582374 438172 582380 438184
rect 454736 438144 582380 438172
rect 454736 438132 454742 438144
rect 582374 438132 582380 438144
rect 582432 438132 582438 438184
rect 360930 431876 360936 431928
rect 360988 431916 360994 431928
rect 580166 431916 580172 431928
rect 360988 431888 580172 431916
rect 360988 431876 360994 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 7558 423620 7564 423632
rect 3384 423592 7564 423620
rect 3384 423580 3390 423592
rect 7558 423580 7564 423592
rect 7616 423580 7622 423632
rect 3326 411204 3332 411256
rect 3384 411244 3390 411256
rect 228542 411244 228548 411256
rect 3384 411216 228548 411244
rect 3384 411204 3390 411216
rect 228542 411204 228548 411216
rect 228600 411204 228606 411256
rect 3326 398760 3332 398812
rect 3384 398800 3390 398812
rect 230014 398800 230020 398812
rect 3384 398772 230020 398800
rect 3384 398760 3390 398772
rect 230014 398760 230020 398772
rect 230072 398760 230078 398812
rect 367738 379448 367744 379500
rect 367796 379488 367802 379500
rect 580166 379488 580172 379500
rect 367796 379460 580172 379488
rect 367796 379448 367802 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3050 372512 3056 372564
rect 3108 372552 3114 372564
rect 229922 372552 229928 372564
rect 3108 372524 229928 372552
rect 3108 372512 3114 372524
rect 229922 372512 229928 372524
rect 229980 372512 229986 372564
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 229830 346372 229836 346384
rect 3384 346344 229836 346372
rect 3384 346332 3390 346344
rect 229830 346332 229836 346344
rect 229888 346332 229894 346384
rect 362218 325592 362224 325644
rect 362276 325632 362282 325644
rect 579890 325632 579896 325644
rect 362276 325604 579896 325632
rect 362276 325592 362282 325604
rect 579890 325592 579896 325604
rect 579948 325592 579954 325644
rect 3326 320084 3332 320136
rect 3384 320124 3390 320136
rect 228450 320124 228456 320136
rect 3384 320096 228456 320124
rect 3384 320084 3390 320096
rect 228450 320084 228456 320096
rect 228508 320084 228514 320136
rect 305362 309136 305368 309188
rect 305420 309176 305426 309188
rect 306190 309176 306196 309188
rect 305420 309148 306196 309176
rect 305420 309136 305426 309148
rect 306190 309136 306196 309148
rect 306248 309136 306254 309188
rect 309134 309136 309140 309188
rect 309192 309176 309198 309188
rect 309410 309176 309416 309188
rect 309192 309148 309416 309176
rect 309192 309136 309198 309148
rect 309410 309136 309416 309148
rect 309468 309136 309474 309188
rect 39298 309068 39304 309120
rect 39356 309108 39362 309120
rect 244458 309108 244464 309120
rect 39356 309080 244464 309108
rect 39356 309068 39362 309080
rect 244458 309068 244464 309080
rect 244516 309068 244522 309120
rect 280062 309068 280068 309120
rect 280120 309108 280126 309120
rect 287606 309108 287612 309120
rect 280120 309080 287612 309108
rect 280120 309068 280126 309080
rect 287606 309068 287612 309080
rect 287664 309068 287670 309120
rect 294966 309068 294972 309120
rect 295024 309108 295030 309120
rect 335814 309108 335820 309120
rect 295024 309080 335820 309108
rect 295024 309068 295030 309080
rect 335814 309068 335820 309080
rect 335872 309068 335878 309120
rect 335998 309068 336004 309120
rect 336056 309108 336062 309120
rect 342346 309108 342352 309120
rect 336056 309080 342352 309108
rect 336056 309068 336062 309080
rect 342346 309068 342352 309080
rect 342404 309068 342410 309120
rect 238018 309000 238024 309052
rect 238076 309040 238082 309052
rect 258258 309040 258264 309052
rect 238076 309012 258264 309040
rect 238076 309000 238082 309012
rect 258258 309000 258264 309012
rect 258316 309000 258322 309052
rect 266446 309000 266452 309052
rect 266504 309040 266510 309052
rect 267458 309040 267464 309052
rect 266504 309012 267464 309040
rect 266504 309000 266510 309012
rect 267458 309000 267464 309012
rect 267516 309000 267522 309052
rect 282638 309000 282644 309052
rect 282696 309040 282702 309052
rect 331858 309040 331864 309052
rect 282696 309012 331864 309040
rect 282696 309000 282702 309012
rect 331858 309000 331864 309012
rect 331916 309000 331922 309052
rect 331950 309000 331956 309052
rect 332008 309040 332014 309052
rect 349890 309040 349896 309052
rect 332008 309012 349896 309040
rect 332008 309000 332014 309012
rect 349890 309000 349896 309012
rect 349948 309000 349954 309052
rect 238202 308932 238208 308984
rect 238260 308972 238266 308984
rect 341794 308972 341800 308984
rect 238260 308944 341800 308972
rect 238260 308932 238266 308944
rect 341794 308932 341800 308944
rect 341852 308932 341858 308984
rect 350626 308972 350632 308984
rect 344986 308944 350632 308972
rect 68278 308864 68284 308916
rect 68336 308904 68342 308916
rect 243170 308904 243176 308916
rect 68336 308876 243176 308904
rect 68336 308864 68342 308876
rect 243170 308864 243176 308876
rect 243228 308864 243234 308916
rect 257982 308864 257988 308916
rect 258040 308904 258046 308916
rect 266446 308904 266452 308916
rect 258040 308876 266452 308904
rect 258040 308864 258046 308876
rect 266446 308864 266452 308876
rect 266504 308864 266510 308916
rect 267090 308864 267096 308916
rect 267148 308904 267154 308916
rect 344986 308904 345014 308944
rect 350626 308932 350632 308944
rect 350684 308932 350690 308984
rect 267148 308876 345014 308904
rect 267148 308864 267154 308876
rect 345842 308864 345848 308916
rect 345900 308904 345906 308916
rect 350166 308904 350172 308916
rect 345900 308876 350172 308904
rect 345900 308864 345906 308876
rect 350166 308864 350172 308876
rect 350224 308864 350230 308916
rect 57238 308796 57244 308848
rect 57296 308836 57302 308848
rect 246666 308836 246672 308848
rect 57296 308808 246672 308836
rect 57296 308796 57302 308808
rect 246666 308796 246672 308808
rect 246724 308796 246730 308848
rect 248138 308796 248144 308848
rect 248196 308836 248202 308848
rect 256050 308836 256056 308848
rect 248196 308808 256056 308836
rect 248196 308796 248202 308808
rect 256050 308796 256056 308808
rect 256108 308796 256114 308848
rect 256142 308796 256148 308848
rect 256200 308836 256206 308848
rect 267274 308836 267280 308848
rect 256200 308808 267280 308836
rect 256200 308796 256206 308808
rect 267274 308796 267280 308808
rect 267332 308796 267338 308848
rect 285030 308796 285036 308848
rect 285088 308836 285094 308848
rect 335998 308836 336004 308848
rect 285088 308808 336004 308836
rect 285088 308796 285094 308808
rect 335998 308796 336004 308808
rect 336056 308796 336062 308848
rect 341058 308836 341064 308848
rect 340846 308808 341064 308836
rect 50338 308728 50344 308780
rect 50396 308768 50402 308780
rect 245562 308768 245568 308780
rect 50396 308740 245568 308768
rect 50396 308728 50402 308740
rect 245562 308728 245568 308740
rect 245620 308728 245626 308780
rect 248414 308728 248420 308780
rect 248472 308768 248478 308780
rect 254946 308768 254952 308780
rect 248472 308740 254952 308768
rect 248472 308728 248478 308740
rect 254946 308728 254952 308740
rect 255004 308728 255010 308780
rect 287606 308728 287612 308780
rect 287664 308768 287670 308780
rect 340846 308768 340874 308808
rect 341058 308796 341064 308808
rect 341116 308796 341122 308848
rect 345290 308796 345296 308848
rect 345348 308836 345354 308848
rect 436830 308836 436836 308848
rect 345348 308808 436836 308836
rect 345348 308796 345354 308808
rect 436830 308796 436836 308808
rect 436888 308796 436894 308848
rect 287664 308740 340874 308768
rect 287664 308728 287670 308740
rect 346394 308728 346400 308780
rect 346452 308768 346458 308780
rect 346452 308740 348004 308768
rect 346452 308728 346458 308740
rect 43438 308660 43444 308712
rect 43496 308700 43502 308712
rect 241698 308700 241704 308712
rect 43496 308672 241704 308700
rect 43496 308660 43502 308672
rect 241698 308660 241704 308672
rect 241756 308660 241762 308712
rect 248046 308660 248052 308712
rect 248104 308700 248110 308712
rect 255498 308700 255504 308712
rect 248104 308672 255504 308700
rect 248104 308660 248110 308672
rect 255498 308660 255504 308672
rect 255556 308660 255562 308712
rect 257430 308660 257436 308712
rect 257488 308700 257494 308712
rect 263962 308700 263968 308712
rect 257488 308672 263968 308700
rect 257488 308660 257494 308672
rect 263962 308660 263968 308672
rect 264020 308660 264026 308712
rect 284110 308660 284116 308712
rect 284168 308700 284174 308712
rect 347130 308700 347136 308712
rect 284168 308672 347136 308700
rect 284168 308660 284174 308672
rect 347130 308660 347136 308672
rect 347188 308660 347194 308712
rect 347976 308700 348004 308740
rect 348050 308728 348056 308780
rect 348108 308768 348114 308780
rect 440602 308768 440608 308780
rect 348108 308740 440608 308768
rect 348108 308728 348114 308740
rect 440602 308728 440608 308740
rect 440660 308728 440666 308780
rect 439590 308700 439596 308712
rect 347976 308672 439596 308700
rect 439590 308660 439596 308672
rect 439648 308660 439654 308712
rect 32398 308592 32404 308644
rect 32456 308632 32462 308644
rect 243722 308632 243728 308644
rect 32456 308604 243728 308632
rect 32456 308592 32462 308604
rect 243722 308592 243728 308604
rect 243780 308592 243786 308644
rect 246666 308592 246672 308644
rect 246724 308632 246730 308644
rect 253842 308632 253848 308644
rect 246724 308604 253848 308632
rect 246724 308592 246730 308604
rect 253842 308592 253848 308604
rect 253900 308592 253906 308644
rect 274542 308592 274548 308644
rect 274600 308632 274606 308644
rect 339954 308632 339960 308644
rect 274600 308604 339960 308632
rect 274600 308592 274606 308604
rect 339954 308592 339960 308604
rect 340012 308592 340018 308644
rect 344094 308592 344100 308644
rect 344152 308632 344158 308644
rect 344922 308632 344928 308644
rect 344152 308604 344928 308632
rect 344152 308592 344158 308604
rect 344922 308592 344928 308604
rect 344980 308592 344986 308644
rect 346486 308592 346492 308644
rect 346544 308632 346550 308644
rect 346946 308632 346952 308644
rect 346544 308604 346952 308632
rect 346544 308592 346550 308604
rect 346946 308592 346952 308604
rect 347004 308592 347010 308644
rect 349246 308592 349252 308644
rect 349304 308632 349310 308644
rect 349522 308632 349528 308644
rect 349304 308604 349528 308632
rect 349304 308592 349310 308604
rect 349522 308592 349528 308604
rect 349580 308592 349586 308644
rect 350166 308592 350172 308644
rect 350224 308632 350230 308644
rect 438118 308632 438124 308644
rect 350224 308604 438124 308632
rect 350224 308592 350230 308604
rect 438118 308592 438124 308604
rect 438176 308592 438182 308644
rect 244918 308524 244924 308576
rect 244976 308564 244982 308576
rect 247034 308564 247040 308576
rect 244976 308536 247040 308564
rect 244976 308524 244982 308536
rect 247034 308524 247040 308536
rect 247092 308524 247098 308576
rect 248322 308564 248328 308576
rect 248156 308536 248328 308564
rect 25498 308456 25504 308508
rect 25556 308496 25562 308508
rect 242986 308496 242992 308508
rect 25556 308468 242992 308496
rect 25556 308456 25562 308468
rect 242986 308456 242992 308468
rect 243044 308456 243050 308508
rect 246574 308456 246580 308508
rect 246632 308496 246638 308508
rect 247218 308496 247224 308508
rect 246632 308468 247224 308496
rect 246632 308456 246638 308468
rect 247218 308456 247224 308468
rect 247276 308456 247282 308508
rect 247586 308456 247592 308508
rect 247644 308456 247650 308508
rect 247770 308456 247776 308508
rect 247828 308456 247834 308508
rect 7558 308388 7564 308440
rect 7616 308428 7622 308440
rect 240778 308428 240784 308440
rect 7616 308400 240784 308428
rect 7616 308388 7622 308400
rect 240778 308388 240784 308400
rect 240836 308388 240842 308440
rect 243078 308388 243084 308440
rect 243136 308428 243142 308440
rect 243538 308428 243544 308440
rect 243136 308400 243544 308428
rect 243136 308388 243142 308400
rect 243538 308388 243544 308400
rect 243596 308388 243602 308440
rect 246298 308388 246304 308440
rect 246356 308388 246362 308440
rect 242986 308320 242992 308372
rect 243044 308360 243050 308372
rect 244090 308360 244096 308372
rect 243044 308332 244096 308360
rect 243044 308320 243050 308332
rect 244090 308320 244096 308332
rect 244148 308320 244154 308372
rect 241606 308252 241612 308304
rect 241664 308292 241670 308304
rect 241790 308292 241796 308304
rect 241664 308264 241796 308292
rect 241664 308252 241670 308264
rect 241790 308252 241796 308264
rect 241848 308252 241854 308304
rect 241974 308252 241980 308304
rect 242032 308292 242038 308304
rect 242434 308292 242440 308304
rect 242032 308264 242440 308292
rect 242032 308252 242038 308264
rect 242434 308252 242440 308264
rect 242492 308252 242498 308304
rect 244550 308252 244556 308304
rect 244608 308292 244614 308304
rect 245378 308292 245384 308304
rect 244608 308264 245384 308292
rect 244608 308252 244614 308264
rect 245378 308252 245384 308264
rect 245436 308252 245442 308304
rect 245930 308252 245936 308304
rect 245988 308292 245994 308304
rect 246316 308292 246344 308388
rect 245988 308264 246344 308292
rect 245988 308252 245994 308264
rect 247218 308252 247224 308304
rect 247276 308292 247282 308304
rect 247604 308292 247632 308456
rect 247276 308264 247632 308292
rect 247276 308252 247282 308264
rect 244458 308184 244464 308236
rect 244516 308224 244522 308236
rect 245194 308224 245200 308236
rect 244516 308196 245200 308224
rect 244516 308184 244522 308196
rect 245194 308184 245200 308196
rect 245252 308184 245258 308236
rect 245838 308184 245844 308236
rect 245896 308224 245902 308236
rect 246850 308224 246856 308236
rect 245896 308196 246856 308224
rect 245896 308184 245902 308196
rect 246850 308184 246856 308196
rect 246908 308184 246914 308236
rect 247402 308184 247408 308236
rect 247460 308224 247466 308236
rect 247788 308224 247816 308456
rect 247954 308252 247960 308304
rect 248012 308292 248018 308304
rect 248156 308292 248184 308536
rect 248322 308524 248328 308536
rect 248380 308524 248386 308576
rect 257154 308564 257160 308576
rect 248616 308536 257160 308564
rect 248414 308496 248420 308508
rect 248012 308264 248184 308292
rect 248248 308468 248420 308496
rect 248012 308252 248018 308264
rect 247460 308196 247816 308224
rect 248248 308224 248276 308468
rect 248414 308456 248420 308468
rect 248472 308456 248478 308508
rect 248322 308388 248328 308440
rect 248380 308428 248386 308440
rect 248616 308428 248644 308536
rect 257154 308524 257160 308536
rect 257212 308524 257218 308576
rect 277118 308524 277124 308576
rect 277176 308564 277182 308576
rect 339402 308564 339408 308576
rect 277176 308536 339408 308564
rect 277176 308524 277182 308536
rect 339402 308524 339408 308536
rect 339460 308524 339466 308576
rect 344186 308524 344192 308576
rect 344244 308564 344250 308576
rect 438026 308564 438032 308576
rect 344244 308536 438032 308564
rect 344244 308524 344250 308536
rect 438026 308524 438032 308536
rect 438084 308524 438090 308576
rect 248782 308456 248788 308508
rect 248840 308496 248846 308508
rect 249058 308496 249064 308508
rect 248840 308468 249064 308496
rect 248840 308456 248846 308468
rect 249058 308456 249064 308468
rect 249116 308456 249122 308508
rect 267826 308456 267832 308508
rect 267884 308496 267890 308508
rect 268194 308496 268200 308508
rect 267884 308468 268200 308496
rect 267884 308456 267890 308468
rect 268194 308456 268200 308468
rect 268252 308456 268258 308508
rect 270494 308456 270500 308508
rect 270552 308496 270558 308508
rect 271506 308496 271512 308508
rect 270552 308468 271512 308496
rect 270552 308456 270558 308468
rect 271506 308456 271512 308468
rect 271564 308456 271570 308508
rect 277302 308456 277308 308508
rect 277360 308496 277366 308508
rect 335998 308496 336004 308508
rect 277360 308468 336004 308496
rect 277360 308456 277366 308468
rect 335998 308456 336004 308468
rect 336056 308456 336062 308508
rect 342346 308456 342352 308508
rect 342404 308496 342410 308508
rect 343266 308496 343272 308508
rect 342404 308468 343272 308496
rect 342404 308456 342410 308468
rect 343266 308456 343272 308468
rect 343324 308456 343330 308508
rect 344738 308456 344744 308508
rect 344796 308496 344802 308508
rect 439498 308496 439504 308508
rect 344796 308468 439504 308496
rect 344796 308456 344802 308468
rect 439498 308456 439504 308468
rect 439556 308456 439562 308508
rect 248380 308400 248644 308428
rect 248380 308388 248386 308400
rect 250254 308388 250260 308440
rect 250312 308428 250318 308440
rect 250898 308428 250904 308440
rect 250312 308400 250904 308428
rect 250312 308388 250318 308400
rect 250898 308388 250904 308400
rect 250956 308388 250962 308440
rect 251174 308388 251180 308440
rect 251232 308428 251238 308440
rect 251818 308428 251824 308440
rect 251232 308400 251824 308428
rect 251232 308388 251238 308400
rect 251818 308388 251824 308400
rect 251876 308388 251882 308440
rect 252646 308388 252652 308440
rect 252704 308428 252710 308440
rect 252922 308428 252928 308440
rect 252704 308400 252928 308428
rect 252704 308388 252710 308400
rect 252922 308388 252928 308400
rect 252980 308388 252986 308440
rect 264606 308388 264612 308440
rect 264664 308428 264670 308440
rect 265066 308428 265072 308440
rect 264664 308400 265072 308428
rect 264664 308388 264670 308400
rect 265066 308388 265072 308400
rect 265124 308388 265130 308440
rect 265158 308388 265164 308440
rect 265216 308428 265222 308440
rect 265434 308428 265440 308440
rect 265216 308400 265440 308428
rect 265216 308388 265222 308400
rect 265434 308388 265440 308400
rect 265492 308388 265498 308440
rect 266446 308388 266452 308440
rect 266504 308428 266510 308440
rect 266906 308428 266912 308440
rect 266504 308400 266912 308428
rect 266504 308388 266510 308400
rect 266906 308388 266912 308400
rect 266964 308388 266970 308440
rect 267734 308388 267740 308440
rect 267792 308428 267798 308440
rect 268746 308428 268752 308440
rect 267792 308400 268752 308428
rect 267792 308388 267798 308400
rect 268746 308388 268752 308400
rect 268804 308388 268810 308440
rect 269298 308388 269304 308440
rect 269356 308428 269362 308440
rect 269850 308428 269856 308440
rect 269356 308400 269856 308428
rect 269356 308388 269362 308400
rect 269850 308388 269856 308400
rect 269908 308388 269914 308440
rect 271230 308388 271236 308440
rect 271288 308428 271294 308440
rect 271874 308428 271880 308440
rect 271288 308400 271880 308428
rect 271288 308388 271294 308400
rect 271874 308388 271880 308400
rect 271932 308388 271938 308440
rect 272150 308388 272156 308440
rect 272208 308428 272214 308440
rect 272978 308428 272984 308440
rect 272208 308400 272984 308428
rect 272208 308388 272214 308400
rect 272978 308388 272984 308400
rect 273036 308388 273042 308440
rect 302326 308388 302332 308440
rect 302384 308428 302390 308440
rect 302602 308428 302608 308440
rect 302384 308400 302608 308428
rect 302384 308388 302390 308400
rect 302602 308388 302608 308400
rect 302660 308388 302666 308440
rect 302694 308388 302700 308440
rect 302752 308428 302758 308440
rect 302970 308428 302976 308440
rect 302752 308400 302976 308428
rect 302752 308388 302758 308400
rect 302970 308388 302976 308400
rect 303028 308388 303034 308440
rect 303798 308388 303804 308440
rect 303856 308428 303862 308440
rect 304810 308428 304816 308440
rect 303856 308400 304816 308428
rect 303856 308388 303862 308400
rect 304810 308388 304816 308400
rect 304868 308388 304874 308440
rect 305270 308388 305276 308440
rect 305328 308428 305334 308440
rect 306098 308428 306104 308440
rect 305328 308400 306104 308428
rect 305328 308388 305334 308400
rect 306098 308388 306104 308400
rect 306156 308388 306162 308440
rect 306190 308388 306196 308440
rect 306248 308428 306254 308440
rect 438854 308428 438860 308440
rect 306248 308400 438860 308428
rect 306248 308388 306254 308400
rect 438854 308388 438860 308400
rect 438912 308388 438918 308440
rect 248414 308320 248420 308372
rect 248472 308360 248478 308372
rect 249610 308360 249616 308372
rect 248472 308332 249616 308360
rect 248472 308320 248478 308332
rect 249610 308320 249616 308332
rect 249668 308320 249674 308372
rect 252830 308320 252836 308372
rect 252888 308360 252894 308372
rect 253474 308360 253480 308372
rect 252888 308332 253480 308360
rect 252888 308320 252894 308332
rect 253474 308320 253480 308332
rect 253532 308320 253538 308372
rect 270678 308320 270684 308372
rect 270736 308360 270742 308372
rect 271322 308360 271328 308372
rect 270736 308332 271328 308360
rect 270736 308320 270742 308332
rect 271322 308320 271328 308332
rect 271380 308320 271386 308372
rect 271966 308320 271972 308372
rect 272024 308360 272030 308372
rect 273162 308360 273168 308372
rect 272024 308332 273168 308360
rect 272024 308320 272030 308332
rect 273162 308320 273168 308332
rect 273220 308320 273226 308372
rect 282822 308320 282828 308372
rect 282880 308360 282886 308372
rect 330938 308360 330944 308372
rect 282880 308332 330944 308360
rect 282880 308320 282886 308332
rect 330938 308320 330944 308332
rect 330996 308320 331002 308372
rect 332502 308320 332508 308372
rect 332560 308360 332566 308372
rect 332560 308332 345014 308360
rect 332560 308320 332566 308332
rect 248598 308252 248604 308304
rect 248656 308292 248662 308304
rect 249242 308292 249248 308304
rect 248656 308264 249248 308292
rect 248656 308252 248662 308264
rect 249242 308252 249248 308264
rect 249300 308252 249306 308304
rect 251450 308252 251456 308304
rect 251508 308292 251514 308304
rect 252186 308292 252192 308304
rect 251508 308264 252192 308292
rect 251508 308252 251514 308264
rect 252186 308252 252192 308264
rect 252244 308252 252250 308304
rect 252554 308252 252560 308304
rect 252612 308292 252618 308304
rect 253106 308292 253112 308304
rect 252612 308264 253112 308292
rect 252612 308252 252618 308264
rect 253106 308252 253112 308264
rect 253164 308252 253170 308304
rect 263594 308252 263600 308304
rect 263652 308292 263658 308304
rect 263962 308292 263968 308304
rect 263652 308264 263968 308292
rect 263652 308252 263658 308264
rect 263962 308252 263968 308264
rect 264020 308252 264026 308304
rect 265066 308252 265072 308304
rect 265124 308292 265130 308304
rect 265986 308292 265992 308304
rect 265124 308264 265992 308292
rect 265124 308252 265130 308264
rect 265986 308252 265992 308264
rect 266044 308252 266050 308304
rect 266354 308252 266360 308304
rect 266412 308292 266418 308304
rect 266906 308292 266912 308304
rect 266412 308264 266912 308292
rect 266412 308252 266418 308264
rect 266906 308252 266912 308264
rect 266964 308252 266970 308304
rect 267918 308252 267924 308304
rect 267976 308292 267982 308304
rect 268286 308292 268292 308304
rect 267976 308264 268292 308292
rect 267976 308252 267982 308264
rect 268286 308252 268292 308264
rect 268344 308252 268350 308304
rect 269114 308252 269120 308304
rect 269172 308292 269178 308304
rect 269574 308292 269580 308304
rect 269172 308264 269580 308292
rect 269172 308252 269178 308264
rect 269574 308252 269580 308264
rect 269632 308252 269638 308304
rect 272242 308252 272248 308304
rect 272300 308292 272306 308304
rect 272426 308292 272432 308304
rect 272300 308264 272432 308292
rect 272300 308252 272306 308264
rect 272426 308252 272432 308264
rect 272484 308252 272490 308304
rect 304994 308252 305000 308304
rect 305052 308292 305058 308304
rect 305546 308292 305552 308304
rect 305052 308264 305552 308292
rect 305052 308252 305058 308264
rect 305546 308252 305552 308264
rect 305604 308252 305610 308304
rect 306558 308252 306564 308304
rect 306616 308292 306622 308304
rect 307202 308292 307208 308304
rect 306616 308264 307208 308292
rect 306616 308252 306622 308264
rect 307202 308252 307208 308264
rect 307260 308252 307266 308304
rect 308214 308252 308220 308304
rect 308272 308292 308278 308304
rect 308674 308292 308680 308304
rect 308272 308264 308680 308292
rect 308272 308252 308278 308264
rect 308674 308252 308680 308264
rect 308732 308252 308738 308304
rect 309134 308252 309140 308304
rect 309192 308292 309198 308304
rect 309962 308292 309968 308304
rect 309192 308264 309968 308292
rect 309192 308252 309198 308264
rect 309962 308252 309968 308264
rect 310020 308252 310026 308304
rect 310698 308252 310704 308304
rect 310756 308292 310762 308304
rect 311710 308292 311716 308304
rect 310756 308264 311716 308292
rect 310756 308252 310762 308264
rect 311710 308252 311716 308264
rect 311768 308252 311774 308304
rect 342530 308252 342536 308304
rect 342588 308292 342594 308304
rect 343082 308292 343088 308304
rect 342588 308264 343088 308292
rect 342588 308252 342594 308264
rect 343082 308252 343088 308264
rect 343140 308252 343146 308304
rect 248248 308196 248368 308224
rect 247460 308184 247466 308196
rect 241790 308116 241796 308168
rect 241848 308156 241854 308168
rect 242802 308156 242808 308168
rect 241848 308128 242808 308156
rect 241848 308116 241854 308128
rect 242802 308116 242808 308128
rect 242860 308116 242866 308168
rect 245654 308116 245660 308168
rect 245712 308156 245718 308168
rect 246206 308156 246212 308168
rect 245712 308128 246212 308156
rect 245712 308116 245718 308128
rect 246206 308116 246212 308128
rect 246264 308116 246270 308168
rect 247310 308116 247316 308168
rect 247368 308156 247374 308168
rect 248230 308156 248236 308168
rect 247368 308128 248236 308156
rect 247368 308116 247374 308128
rect 248230 308116 248236 308128
rect 248288 308116 248294 308168
rect 243630 308048 243636 308100
rect 243688 308088 243694 308100
rect 248340 308088 248368 308196
rect 252922 308184 252928 308236
rect 252980 308224 252986 308236
rect 253658 308224 253664 308236
rect 252980 308196 253664 308224
rect 252980 308184 252986 308196
rect 253658 308184 253664 308196
rect 253716 308184 253722 308236
rect 263778 308184 263784 308236
rect 263836 308224 263842 308236
rect 264698 308224 264704 308236
rect 263836 308196 264704 308224
rect 263836 308184 263842 308196
rect 264698 308184 264704 308196
rect 264756 308184 264762 308236
rect 268378 308184 268384 308236
rect 268436 308224 268442 308236
rect 272794 308224 272800 308236
rect 268436 308196 272800 308224
rect 268436 308184 268442 308196
rect 272794 308184 272800 308196
rect 272852 308184 272858 308236
rect 302206 308196 316724 308224
rect 265434 308116 265440 308168
rect 265492 308156 265498 308168
rect 266170 308156 266176 308168
rect 265492 308128 266176 308156
rect 265492 308116 265498 308128
rect 266170 308116 266176 308128
rect 266228 308116 266234 308168
rect 266630 308116 266636 308168
rect 266688 308156 266694 308168
rect 266998 308156 267004 308168
rect 266688 308128 267004 308156
rect 266688 308116 266694 308128
rect 266998 308116 267004 308128
rect 267056 308116 267062 308168
rect 267918 308116 267924 308168
rect 267976 308156 267982 308168
rect 268562 308156 268568 308168
rect 267976 308128 268568 308156
rect 267976 308116 267982 308128
rect 268562 308116 268568 308128
rect 268620 308116 268626 308168
rect 269390 308116 269396 308168
rect 269448 308156 269454 308168
rect 269942 308156 269948 308168
rect 269448 308128 269948 308156
rect 269448 308116 269454 308128
rect 269942 308116 269948 308128
rect 270000 308116 270006 308168
rect 272242 308116 272248 308168
rect 272300 308156 272306 308168
rect 272610 308156 272616 308168
rect 272300 308128 272616 308156
rect 272300 308116 272306 308128
rect 272610 308116 272616 308128
rect 272668 308116 272674 308168
rect 250162 308088 250168 308100
rect 243688 308060 248368 308088
rect 249812 308060 250168 308088
rect 243688 308048 243694 308060
rect 249812 308032 249840 308060
rect 250162 308048 250168 308060
rect 250220 308048 250226 308100
rect 253198 308048 253204 308100
rect 253256 308088 253262 308100
rect 258626 308088 258632 308100
rect 253256 308060 258632 308088
rect 253256 308048 253262 308060
rect 258626 308048 258632 308060
rect 258684 308048 258690 308100
rect 266538 308048 266544 308100
rect 266596 308088 266602 308100
rect 267642 308088 267648 308100
rect 266596 308060 267648 308088
rect 266596 308048 266602 308060
rect 267642 308048 267648 308060
rect 267700 308048 267706 308100
rect 286042 308048 286048 308100
rect 286100 308088 286106 308100
rect 291838 308088 291844 308100
rect 286100 308060 291844 308088
rect 286100 308048 286106 308060
rect 291838 308048 291844 308060
rect 291896 308048 291902 308100
rect 291930 308048 291936 308100
rect 291988 308088 291994 308100
rect 293494 308088 293500 308100
rect 291988 308060 293500 308088
rect 291988 308048 291994 308060
rect 293494 308048 293500 308060
rect 293552 308048 293558 308100
rect 240502 307980 240508 308032
rect 240560 308020 240566 308032
rect 241330 308020 241336 308032
rect 240560 307992 241336 308020
rect 240560 307980 240566 307992
rect 241330 307980 241336 307992
rect 241388 307980 241394 308032
rect 243722 307980 243728 308032
rect 243780 308020 243786 308032
rect 245010 308020 245016 308032
rect 243780 307992 245016 308020
rect 243780 307980 243786 307992
rect 245010 307980 245016 307992
rect 245068 307980 245074 308032
rect 248874 307980 248880 308032
rect 248932 308020 248938 308032
rect 249426 308020 249432 308032
rect 248932 307992 249432 308020
rect 248932 307980 248938 307992
rect 249426 307980 249432 307992
rect 249484 307980 249490 308032
rect 249794 307980 249800 308032
rect 249852 307980 249858 308032
rect 249886 307980 249892 308032
rect 249944 308020 249950 308032
rect 250530 308020 250536 308032
rect 249944 307992 250536 308020
rect 249944 307980 249950 307992
rect 250530 307980 250536 307992
rect 250588 307980 250594 308032
rect 265250 307980 265256 308032
rect 265308 308020 265314 308032
rect 265802 308020 265808 308032
rect 265308 307992 265808 308020
rect 265308 307980 265314 307992
rect 265802 307980 265808 307992
rect 265860 307980 265866 308032
rect 269390 307980 269396 308032
rect 269448 308020 269454 308032
rect 270218 308020 270224 308032
rect 269448 307992 270224 308020
rect 269448 307980 269454 307992
rect 270218 307980 270224 307992
rect 270276 307980 270282 308032
rect 280706 308020 280712 308032
rect 273226 307992 280712 308020
rect 242158 307912 242164 307964
rect 242216 307952 242222 307964
rect 248322 307952 248328 307964
rect 242216 307924 248328 307952
rect 242216 307912 242222 307924
rect 248322 307912 248328 307924
rect 248380 307912 248386 307964
rect 250162 307912 250168 307964
rect 250220 307952 250226 307964
rect 250714 307952 250720 307964
rect 250220 307924 250720 307952
rect 250220 307912 250226 307924
rect 250714 307912 250720 307924
rect 250772 307912 250778 307964
rect 254670 307844 254676 307896
rect 254728 307884 254734 307896
rect 258442 307884 258448 307896
rect 254728 307856 258448 307884
rect 254728 307844 254734 307856
rect 258442 307844 258448 307856
rect 258500 307844 258506 307896
rect 246298 307776 246304 307828
rect 246356 307816 246362 307828
rect 246666 307816 246672 307828
rect 246356 307788 246672 307816
rect 246356 307776 246362 307788
rect 246666 307776 246672 307788
rect 246724 307776 246730 307828
rect 247678 307776 247684 307828
rect 247736 307816 247742 307828
rect 248138 307816 248144 307828
rect 247736 307788 248144 307816
rect 247736 307776 247742 307788
rect 248138 307776 248144 307788
rect 248196 307776 248202 307828
rect 255958 307776 255964 307828
rect 256016 307816 256022 307828
rect 256970 307816 256976 307828
rect 256016 307788 256976 307816
rect 256016 307776 256022 307788
rect 256970 307776 256976 307788
rect 257028 307776 257034 307828
rect 260190 307776 260196 307828
rect 260248 307816 260254 307828
rect 262306 307816 262312 307828
rect 260248 307788 262312 307816
rect 260248 307776 260254 307788
rect 262306 307776 262312 307788
rect 262364 307776 262370 307828
rect 265618 307776 265624 307828
rect 265676 307816 265682 307828
rect 269206 307816 269212 307828
rect 265676 307788 269212 307816
rect 265676 307776 265682 307788
rect 269206 307776 269212 307788
rect 269264 307776 269270 307828
rect 269758 307776 269764 307828
rect 269816 307816 269822 307828
rect 273226 307816 273254 307992
rect 280706 307980 280712 307992
rect 280764 307980 280770 308032
rect 290734 307980 290740 308032
rect 290792 308020 290798 308032
rect 302206 308020 302234 308196
rect 305086 308116 305092 308168
rect 305144 308156 305150 308168
rect 305914 308156 305920 308168
rect 305144 308128 305920 308156
rect 305144 308116 305150 308128
rect 305914 308116 305920 308128
rect 305972 308116 305978 308168
rect 306650 308116 306656 308168
rect 306708 308156 306714 308168
rect 307018 308156 307024 308168
rect 306708 308128 307024 308156
rect 306708 308116 306714 308128
rect 307018 308116 307024 308128
rect 307076 308116 307082 308168
rect 308030 308116 308036 308168
rect 308088 308156 308094 308168
rect 308398 308156 308404 308168
rect 308088 308128 308404 308156
rect 308088 308116 308094 308128
rect 308398 308116 308404 308128
rect 308456 308116 308462 308168
rect 309318 308116 309324 308168
rect 309376 308156 309382 308168
rect 310330 308156 310336 308168
rect 309376 308128 310336 308156
rect 309376 308116 309382 308128
rect 310330 308116 310336 308128
rect 310388 308116 310394 308168
rect 306374 308048 306380 308100
rect 306432 308088 306438 308100
rect 307570 308088 307576 308100
rect 306432 308060 307576 308088
rect 306432 308048 306438 308060
rect 307570 308048 307576 308060
rect 307628 308048 307634 308100
rect 307846 308048 307852 308100
rect 307904 308088 307910 308100
rect 309042 308088 309048 308100
rect 307904 308060 309048 308088
rect 307904 308048 307910 308060
rect 309042 308048 309048 308060
rect 309100 308048 309106 308100
rect 290792 307992 302234 308020
rect 290792 307980 290798 307992
rect 304074 307980 304080 308032
rect 304132 308020 304138 308032
rect 304626 308020 304632 308032
rect 304132 307992 304632 308020
rect 304132 307980 304138 307992
rect 304626 307980 304632 307992
rect 304684 307980 304690 308032
rect 307754 307980 307760 308032
rect 307812 308020 307818 308032
rect 308858 308020 308864 308032
rect 307812 307992 308864 308020
rect 307812 307980 307818 307992
rect 308858 307980 308864 307992
rect 308916 307980 308922 308032
rect 310606 307980 310612 308032
rect 310664 308020 310670 308032
rect 311066 308020 311072 308032
rect 310664 307992 311072 308020
rect 310664 307980 310670 307992
rect 311066 307980 311072 307992
rect 311124 307980 311130 308032
rect 311710 307980 311716 308032
rect 311768 308020 311774 308032
rect 312446 308020 312452 308032
rect 311768 307992 312452 308020
rect 311768 307980 311774 307992
rect 312446 307980 312452 307992
rect 312504 307980 312510 308032
rect 286226 307912 286232 307964
rect 286284 307952 286290 307964
rect 293310 307952 293316 307964
rect 286284 307924 293316 307952
rect 286284 307912 286290 307924
rect 293310 307912 293316 307924
rect 293368 307912 293374 307964
rect 295426 307912 295432 307964
rect 295484 307952 295490 307964
rect 297266 307952 297272 307964
rect 295484 307924 297272 307952
rect 295484 307912 295490 307924
rect 297266 307912 297272 307924
rect 297324 307912 297330 307964
rect 302786 307912 302792 307964
rect 302844 307952 302850 307964
rect 303522 307952 303528 307964
rect 302844 307924 303528 307952
rect 302844 307912 302850 307924
rect 303522 307912 303528 307924
rect 303580 307912 303586 307964
rect 303890 307912 303896 307964
rect 303948 307952 303954 307964
rect 304442 307952 304448 307964
rect 303948 307924 304448 307952
rect 303948 307912 303954 307924
rect 304442 307912 304448 307924
rect 304500 307912 304506 307964
rect 310698 307912 310704 307964
rect 310756 307952 310762 307964
rect 311434 307952 311440 307964
rect 310756 307924 311440 307952
rect 310756 307912 310762 307924
rect 311434 307912 311440 307924
rect 311492 307912 311498 307964
rect 278222 307844 278228 307896
rect 278280 307884 278286 307896
rect 279786 307884 279792 307896
rect 278280 307856 279792 307884
rect 278280 307844 278286 307856
rect 279786 307844 279792 307856
rect 279844 307844 279850 307896
rect 279878 307844 279884 307896
rect 279936 307884 279942 307896
rect 281258 307884 281264 307896
rect 279936 307856 281264 307884
rect 279936 307844 279942 307856
rect 281258 307844 281264 307856
rect 281316 307844 281322 307896
rect 285122 307844 285128 307896
rect 285180 307884 285186 307896
rect 287790 307884 287796 307896
rect 285180 307856 287796 307884
rect 285180 307844 285186 307856
rect 287790 307844 287796 307856
rect 287848 307844 287854 307896
rect 294690 307844 294696 307896
rect 294748 307884 294754 307896
rect 296254 307884 296260 307896
rect 294748 307856 296260 307884
rect 294748 307844 294754 307856
rect 296254 307844 296260 307856
rect 296312 307844 296318 307896
rect 302602 307844 302608 307896
rect 302660 307884 302666 307896
rect 303338 307884 303344 307896
rect 302660 307856 303344 307884
rect 302660 307844 302666 307856
rect 303338 307844 303344 307856
rect 303396 307844 303402 307896
rect 303706 307844 303712 307896
rect 303764 307884 303770 307896
rect 304258 307884 304264 307896
rect 303764 307856 304264 307884
rect 303764 307844 303770 307856
rect 304258 307844 304264 307856
rect 304316 307844 304322 307896
rect 310790 307844 310796 307896
rect 310848 307884 310854 307896
rect 311802 307884 311808 307896
rect 310848 307856 311808 307884
rect 310848 307844 310854 307856
rect 311802 307844 311808 307856
rect 311860 307844 311866 307896
rect 316696 307884 316724 308196
rect 321462 308184 321468 308236
rect 321520 308224 321526 308236
rect 321830 308224 321836 308236
rect 321520 308196 321836 308224
rect 321520 308184 321526 308196
rect 321830 308184 321836 308196
rect 321888 308184 321894 308236
rect 335814 308184 335820 308236
rect 335872 308224 335878 308236
rect 343450 308224 343456 308236
rect 335872 308196 343456 308224
rect 335872 308184 335878 308196
rect 343450 308184 343456 308196
rect 343508 308184 343514 308236
rect 341426 308116 341432 308168
rect 341484 308156 341490 308168
rect 342162 308156 342168 308168
rect 341484 308128 342168 308156
rect 341484 308116 341490 308128
rect 342162 308116 342168 308128
rect 342220 308116 342226 308168
rect 344986 308156 345014 308332
rect 345198 308320 345204 308372
rect 345256 308360 345262 308372
rect 345658 308360 345664 308372
rect 345256 308332 345664 308360
rect 345256 308320 345262 308332
rect 345658 308320 345664 308332
rect 345716 308320 345722 308372
rect 346946 308320 346952 308372
rect 347004 308360 347010 308372
rect 347682 308360 347688 308372
rect 347004 308332 347688 308360
rect 347004 308320 347010 308332
rect 347682 308320 347688 308332
rect 347740 308320 347746 308372
rect 348050 308320 348056 308372
rect 348108 308360 348114 308372
rect 348418 308360 348424 308372
rect 348108 308332 348424 308360
rect 348108 308320 348114 308332
rect 348418 308320 348424 308332
rect 348476 308320 348482 308372
rect 349154 308320 349160 308372
rect 349212 308360 349218 308372
rect 349614 308360 349620 308372
rect 349212 308332 349620 308360
rect 349212 308320 349218 308332
rect 349614 308320 349620 308332
rect 349672 308320 349678 308372
rect 345106 308252 345112 308304
rect 345164 308292 345170 308304
rect 346210 308292 346216 308304
rect 345164 308264 346216 308292
rect 345164 308252 345170 308264
rect 346210 308252 346216 308264
rect 346268 308252 346274 308304
rect 346670 308252 346676 308304
rect 346728 308292 346734 308304
rect 347498 308292 347504 308304
rect 346728 308264 347504 308292
rect 346728 308252 346734 308264
rect 347498 308252 347504 308264
rect 347556 308252 347562 308304
rect 348234 308252 348240 308304
rect 348292 308292 348298 308304
rect 348786 308292 348792 308304
rect 348292 308264 348792 308292
rect 348292 308252 348298 308264
rect 348786 308252 348792 308264
rect 348844 308252 348850 308304
rect 349338 308252 349344 308304
rect 349396 308292 349402 308304
rect 349706 308292 349712 308304
rect 349396 308264 349712 308292
rect 349396 308252 349402 308264
rect 349706 308252 349712 308264
rect 349764 308252 349770 308304
rect 349430 308184 349436 308236
rect 349488 308224 349494 308236
rect 350258 308224 350264 308236
rect 349488 308196 350264 308224
rect 349488 308184 349494 308196
rect 350258 308184 350264 308196
rect 350316 308184 350322 308236
rect 350442 308156 350448 308168
rect 344986 308128 350448 308156
rect 350442 308116 350448 308128
rect 350500 308116 350506 308168
rect 341242 308048 341248 308100
rect 341300 308088 341306 308100
rect 341978 308088 341984 308100
rect 341300 308060 341984 308088
rect 341300 308048 341306 308060
rect 341978 308048 341984 308060
rect 342036 308048 342042 308100
rect 316862 307912 316868 307964
rect 316920 307952 316926 307964
rect 343634 307952 343640 307964
rect 316920 307924 343640 307952
rect 316920 307912 316926 307924
rect 343634 307912 343640 307924
rect 343692 307912 343698 307964
rect 331122 307884 331128 307896
rect 316696 307856 331128 307884
rect 331122 307844 331128 307856
rect 331180 307844 331186 307896
rect 269816 307788 273254 307816
rect 269816 307776 269822 307788
rect 273990 307776 273996 307828
rect 274048 307816 274054 307828
rect 275002 307816 275008 307828
rect 274048 307788 275008 307816
rect 274048 307776 274054 307788
rect 275002 307776 275008 307788
rect 275060 307776 275066 307828
rect 275462 307776 275468 307828
rect 275520 307816 275526 307828
rect 276106 307816 276112 307828
rect 275520 307788 276112 307816
rect 275520 307776 275526 307788
rect 276106 307776 276112 307788
rect 276164 307776 276170 307828
rect 279694 307776 279700 307828
rect 279752 307816 279758 307828
rect 280338 307816 280344 307828
rect 279752 307788 280344 307816
rect 279752 307776 279758 307788
rect 280338 307776 280344 307788
rect 280396 307776 280402 307828
rect 280982 307776 280988 307828
rect 281040 307816 281046 307828
rect 282730 307816 282736 307828
rect 281040 307788 282736 307816
rect 281040 307776 281046 307788
rect 282730 307776 282736 307788
rect 282788 307776 282794 307828
rect 284202 307776 284208 307828
rect 284260 307816 284266 307828
rect 284478 307816 284484 307828
rect 284260 307788 284484 307816
rect 284260 307776 284266 307788
rect 284478 307776 284484 307788
rect 284536 307776 284542 307828
rect 285306 307776 285312 307828
rect 285364 307816 285370 307828
rect 286318 307816 286324 307828
rect 285364 307788 286324 307816
rect 285364 307776 285370 307788
rect 286318 307776 286324 307788
rect 286376 307776 286382 307828
rect 288802 307776 288808 307828
rect 288860 307816 288866 307828
rect 291930 307816 291936 307828
rect 288860 307788 291936 307816
rect 288860 307776 288866 307788
rect 291930 307776 291936 307788
rect 291988 307776 291994 307828
rect 293586 307776 293592 307828
rect 293644 307816 293650 307828
rect 294598 307816 294604 307828
rect 293644 307788 294604 307816
rect 293644 307776 293650 307788
rect 294598 307776 294604 307788
rect 294656 307776 294662 307828
rect 295242 307776 295248 307828
rect 295300 307816 295306 307828
rect 296070 307816 296076 307828
rect 295300 307788 296076 307816
rect 295300 307776 295306 307788
rect 296070 307776 296076 307788
rect 296128 307776 296134 307828
rect 302418 307776 302424 307828
rect 302476 307816 302482 307828
rect 303154 307816 303160 307828
rect 302476 307788 303160 307816
rect 302476 307776 302482 307788
rect 303154 307776 303160 307788
rect 303212 307776 303218 307828
rect 310514 307776 310520 307828
rect 310572 307816 310578 307828
rect 311618 307816 311624 307828
rect 310572 307788 311624 307816
rect 310572 307776 310578 307788
rect 311618 307776 311624 307788
rect 311676 307776 311682 307828
rect 312906 307776 312912 307828
rect 312964 307816 312970 307828
rect 315298 307816 315304 307828
rect 312964 307788 315304 307816
rect 312964 307776 312970 307788
rect 315298 307776 315304 307788
rect 315356 307776 315362 307828
rect 335998 307776 336004 307828
rect 336056 307816 336062 307828
rect 344370 307816 344376 307828
rect 336056 307788 344376 307816
rect 336056 307776 336062 307788
rect 344370 307776 344376 307788
rect 344428 307776 344434 307828
rect 269206 307640 269212 307692
rect 269264 307680 269270 307692
rect 270402 307680 270408 307692
rect 269264 307652 270408 307680
rect 269264 307640 269270 307652
rect 270402 307640 270408 307652
rect 270460 307640 270466 307692
rect 270586 307368 270592 307420
rect 270644 307408 270650 307420
rect 270954 307408 270960 307420
rect 270644 307380 270960 307408
rect 270644 307368 270650 307380
rect 270954 307368 270960 307380
rect 271012 307368 271018 307420
rect 64874 307232 64880 307284
rect 64932 307272 64938 307284
rect 249794 307272 249800 307284
rect 64932 307244 249800 307272
rect 64932 307232 64938 307244
rect 249794 307232 249800 307244
rect 249852 307232 249858 307284
rect 52454 307164 52460 307216
rect 52512 307204 52518 307216
rect 247954 307204 247960 307216
rect 52512 307176 247960 307204
rect 52512 307164 52518 307176
rect 247954 307164 247960 307176
rect 248012 307164 248018 307216
rect 31018 307096 31024 307148
rect 31076 307136 31082 307148
rect 244734 307136 244740 307148
rect 31076 307108 244740 307136
rect 31076 307096 31082 307108
rect 244734 307096 244740 307108
rect 244792 307096 244798 307148
rect 314746 307096 314752 307148
rect 314804 307136 314810 307148
rect 478138 307136 478144 307148
rect 314804 307108 478144 307136
rect 314804 307096 314810 307108
rect 478138 307096 478144 307108
rect 478196 307096 478202 307148
rect 8938 307028 8944 307080
rect 8996 307068 9002 307080
rect 240134 307068 240140 307080
rect 8996 307040 240140 307068
rect 8996 307028 9002 307040
rect 240134 307028 240140 307040
rect 240192 307028 240198 307080
rect 316218 307028 316224 307080
rect 316276 307068 316282 307080
rect 489914 307068 489920 307080
rect 316276 307040 489920 307068
rect 316276 307028 316282 307040
rect 489914 307028 489920 307040
rect 489972 307028 489978 307080
rect 253934 306960 253940 307012
rect 253992 307000 253998 307012
rect 254210 307000 254216 307012
rect 253992 306972 254216 307000
rect 253992 306960 253998 306972
rect 254210 306960 254216 306972
rect 254268 306960 254274 307012
rect 277762 307000 277768 307012
rect 277688 306972 277768 307000
rect 251542 306824 251548 306876
rect 251600 306864 251606 306876
rect 252370 306864 252376 306876
rect 251600 306836 252376 306864
rect 251600 306824 251606 306836
rect 252370 306824 252376 306836
rect 252428 306824 252434 306876
rect 277688 306808 277716 306972
rect 277762 306960 277768 306972
rect 277820 306960 277826 307012
rect 319070 306824 319076 306876
rect 319128 306864 319134 306876
rect 319346 306864 319352 306876
rect 319128 306836 319352 306864
rect 319128 306824 319134 306836
rect 319346 306824 319352 306836
rect 319404 306824 319410 306876
rect 270954 306756 270960 306808
rect 271012 306796 271018 306808
rect 271690 306796 271696 306808
rect 271012 306768 271696 306796
rect 271012 306756 271018 306768
rect 271690 306756 271696 306768
rect 271748 306756 271754 306808
rect 277670 306756 277676 306808
rect 277728 306756 277734 306808
rect 299842 306688 299848 306740
rect 299900 306688 299906 306740
rect 258810 306552 258816 306604
rect 258868 306552 258874 306604
rect 268102 306552 268108 306604
rect 268160 306592 268166 306604
rect 268930 306592 268936 306604
rect 268160 306564 268936 306592
rect 268160 306552 268166 306564
rect 268930 306552 268936 306564
rect 268988 306552 268994 306604
rect 296714 306552 296720 306604
rect 296772 306592 296778 306604
rect 297174 306592 297180 306604
rect 296772 306564 297180 306592
rect 296772 306552 296778 306564
rect 297174 306552 297180 306564
rect 297232 306552 297238 306604
rect 255498 306348 255504 306400
rect 255556 306388 255562 306400
rect 255866 306388 255872 306400
rect 255556 306360 255872 306388
rect 255556 306348 255562 306360
rect 255866 306348 255872 306360
rect 255924 306348 255930 306400
rect 258258 306348 258264 306400
rect 258316 306388 258322 306400
rect 258828 306388 258856 306552
rect 277578 306484 277584 306536
rect 277636 306524 277642 306536
rect 277854 306524 277860 306536
rect 277636 306496 277860 306524
rect 277636 306484 277642 306496
rect 277854 306484 277860 306496
rect 277912 306484 277918 306536
rect 285674 306484 285680 306536
rect 285732 306524 285738 306536
rect 286042 306524 286048 306536
rect 285732 306496 286048 306524
rect 285732 306484 285738 306496
rect 286042 306484 286048 306496
rect 286100 306484 286106 306536
rect 286134 306484 286140 306536
rect 286192 306524 286198 306536
rect 286594 306524 286600 306536
rect 286192 306496 286600 306524
rect 286192 306484 286198 306496
rect 286594 306484 286600 306496
rect 286652 306484 286658 306536
rect 289814 306484 289820 306536
rect 289872 306524 289878 306536
rect 291010 306524 291016 306536
rect 289872 306496 291016 306524
rect 289872 306484 289878 306496
rect 291010 306484 291016 306496
rect 291068 306484 291074 306536
rect 292942 306484 292948 306536
rect 293000 306524 293006 306536
rect 293218 306524 293224 306536
rect 293000 306496 293224 306524
rect 293000 306484 293006 306496
rect 293218 306484 293224 306496
rect 293276 306484 293282 306536
rect 299860 306468 299888 306688
rect 329374 306552 329380 306604
rect 329432 306592 329438 306604
rect 332962 306592 332968 306604
rect 329432 306564 332968 306592
rect 329432 306552 329438 306564
rect 332962 306552 332968 306564
rect 333020 306552 333026 306604
rect 314746 306484 314752 306536
rect 314804 306524 314810 306536
rect 315666 306524 315672 306536
rect 314804 306496 315672 306524
rect 314804 306484 314810 306496
rect 315666 306484 315672 306496
rect 315724 306484 315730 306536
rect 317506 306484 317512 306536
rect 317564 306524 317570 306536
rect 317966 306524 317972 306536
rect 317564 306496 317972 306524
rect 317564 306484 317570 306496
rect 317966 306484 317972 306496
rect 318024 306484 318030 306536
rect 328454 306484 328460 306536
rect 328512 306524 328518 306536
rect 329466 306524 329472 306536
rect 328512 306496 329472 306524
rect 328512 306484 328518 306496
rect 329466 306484 329472 306496
rect 329524 306484 329530 306536
rect 259546 306416 259552 306468
rect 259604 306456 259610 306468
rect 259914 306456 259920 306468
rect 259604 306428 259920 306456
rect 259604 306416 259610 306428
rect 259914 306416 259920 306428
rect 259972 306416 259978 306468
rect 277486 306416 277492 306468
rect 277544 306456 277550 306468
rect 278130 306456 278136 306468
rect 277544 306428 278136 306456
rect 277544 306416 277550 306428
rect 278130 306416 278136 306428
rect 278188 306416 278194 306468
rect 278958 306416 278964 306468
rect 279016 306456 279022 306468
rect 279234 306456 279240 306468
rect 279016 306428 279240 306456
rect 279016 306416 279022 306428
rect 279234 306416 279240 306428
rect 279292 306416 279298 306468
rect 286410 306456 286416 306468
rect 285692 306428 286416 306456
rect 285692 306400 285720 306428
rect 286410 306416 286416 306428
rect 286468 306416 286474 306468
rect 289906 306416 289912 306468
rect 289964 306456 289970 306468
rect 290366 306456 290372 306468
rect 289964 306428 290372 306456
rect 289964 306416 289970 306428
rect 290366 306416 290372 306428
rect 290424 306416 290430 306468
rect 291194 306416 291200 306468
rect 291252 306456 291258 306468
rect 291470 306456 291476 306468
rect 291252 306428 291476 306456
rect 291252 306416 291258 306428
rect 291470 306416 291476 306428
rect 291528 306416 291534 306468
rect 292666 306416 292672 306468
rect 292724 306456 292730 306468
rect 293402 306456 293408 306468
rect 292724 306428 293408 306456
rect 292724 306416 292730 306428
rect 293402 306416 293408 306428
rect 293460 306416 293466 306468
rect 293954 306416 293960 306468
rect 294012 306456 294018 306468
rect 295886 306456 295892 306468
rect 294012 306428 295892 306456
rect 294012 306416 294018 306428
rect 295886 306416 295892 306428
rect 295944 306416 295950 306468
rect 298186 306416 298192 306468
rect 298244 306456 298250 306468
rect 298462 306456 298468 306468
rect 298244 306428 298468 306456
rect 298244 306416 298250 306428
rect 298462 306416 298468 306428
rect 298520 306416 298526 306468
rect 299842 306416 299848 306468
rect 299900 306416 299906 306468
rect 300854 306416 300860 306468
rect 300912 306456 300918 306468
rect 302050 306456 302056 306468
rect 300912 306428 302056 306456
rect 300912 306416 300918 306428
rect 302050 306416 302056 306428
rect 302108 306416 302114 306468
rect 314838 306416 314844 306468
rect 314896 306456 314902 306468
rect 315482 306456 315488 306468
rect 314896 306428 315488 306456
rect 314896 306416 314902 306428
rect 315482 306416 315488 306428
rect 315540 306416 315546 306468
rect 316218 306416 316224 306468
rect 316276 306456 316282 306468
rect 316586 306456 316592 306468
rect 316276 306428 316592 306456
rect 316276 306416 316282 306428
rect 316586 306416 316592 306428
rect 316644 306416 316650 306468
rect 320266 306416 320272 306468
rect 320324 306456 320330 306468
rect 320726 306456 320732 306468
rect 320324 306428 320732 306456
rect 320324 306416 320330 306428
rect 320726 306416 320732 306428
rect 320784 306416 320790 306468
rect 321738 306416 321744 306468
rect 321796 306456 321802 306468
rect 322198 306456 322204 306468
rect 321796 306428 322204 306456
rect 321796 306416 321802 306428
rect 322198 306416 322204 306428
rect 322256 306416 322262 306468
rect 324498 306416 324504 306468
rect 324556 306456 324562 306468
rect 325142 306456 325148 306468
rect 324556 306428 325148 306456
rect 324556 306416 324562 306428
rect 325142 306416 325148 306428
rect 325200 306416 325206 306468
rect 325878 306416 325884 306468
rect 325936 306456 325942 306468
rect 326338 306456 326344 306468
rect 325936 306428 326344 306456
rect 325936 306416 325942 306428
rect 326338 306416 326344 306428
rect 326396 306416 326402 306468
rect 327442 306416 327448 306468
rect 327500 306456 327506 306468
rect 328086 306456 328092 306468
rect 327500 306428 328092 306456
rect 327500 306416 327506 306428
rect 328086 306416 328092 306428
rect 328144 306416 328150 306468
rect 328546 306416 328552 306468
rect 328604 306456 328610 306468
rect 329006 306456 329012 306468
rect 328604 306428 329012 306456
rect 328604 306416 328610 306428
rect 329006 306416 329012 306428
rect 329064 306416 329070 306468
rect 332686 306416 332692 306468
rect 332744 306456 332750 306468
rect 333698 306456 333704 306468
rect 332744 306428 333704 306456
rect 332744 306416 332750 306428
rect 333698 306416 333704 306428
rect 333756 306416 333762 306468
rect 334342 306416 334348 306468
rect 334400 306456 334406 306468
rect 334618 306456 334624 306468
rect 334400 306428 334624 306456
rect 334400 306416 334406 306428
rect 334618 306416 334624 306428
rect 334676 306416 334682 306468
rect 348602 306456 348608 306468
rect 347976 306428 348608 306456
rect 347976 306400 348004 306428
rect 348602 306416 348608 306428
rect 348660 306416 348666 306468
rect 258316 306360 258856 306388
rect 258316 306348 258322 306360
rect 259454 306348 259460 306400
rect 259512 306388 259518 306400
rect 260466 306388 260472 306400
rect 259512 306360 260472 306388
rect 259512 306348 259518 306360
rect 260466 306348 260472 306360
rect 260524 306348 260530 306400
rect 261110 306348 261116 306400
rect 261168 306388 261174 306400
rect 261938 306388 261944 306400
rect 261168 306360 261944 306388
rect 261168 306348 261174 306360
rect 261938 306348 261944 306360
rect 261996 306348 262002 306400
rect 262306 306348 262312 306400
rect 262364 306388 262370 306400
rect 263042 306388 263048 306400
rect 262364 306360 263048 306388
rect 262364 306348 262370 306360
rect 263042 306348 263048 306360
rect 263100 306348 263106 306400
rect 273254 306348 273260 306400
rect 273312 306388 273318 306400
rect 274266 306388 274272 306400
rect 273312 306360 274272 306388
rect 273312 306348 273318 306360
rect 274266 306348 274272 306360
rect 274324 306348 274330 306400
rect 274726 306348 274732 306400
rect 274784 306388 274790 306400
rect 275922 306388 275928 306400
rect 274784 306360 275928 306388
rect 274784 306348 274790 306360
rect 275922 306348 275928 306360
rect 275980 306348 275986 306400
rect 276198 306348 276204 306400
rect 276256 306388 276262 306400
rect 277210 306388 277216 306400
rect 276256 306360 277216 306388
rect 276256 306348 276262 306360
rect 277210 306348 277216 306360
rect 277268 306348 277274 306400
rect 281718 306348 281724 306400
rect 281776 306388 281782 306400
rect 282362 306388 282368 306400
rect 281776 306360 282368 306388
rect 281776 306348 281782 306360
rect 282362 306348 282368 306360
rect 282420 306348 282426 306400
rect 284662 306348 284668 306400
rect 284720 306388 284726 306400
rect 285490 306388 285496 306400
rect 284720 306360 285496 306388
rect 284720 306348 284726 306360
rect 285490 306348 285496 306360
rect 285548 306348 285554 306400
rect 285674 306348 285680 306400
rect 285732 306348 285738 306400
rect 285950 306348 285956 306400
rect 286008 306388 286014 306400
rect 286778 306388 286784 306400
rect 286008 306360 286784 306388
rect 286008 306348 286014 306360
rect 286778 306348 286784 306360
rect 286836 306348 286842 306400
rect 287054 306348 287060 306400
rect 287112 306388 287118 306400
rect 287882 306388 287888 306400
rect 287112 306360 287888 306388
rect 287112 306348 287118 306360
rect 287882 306348 287888 306360
rect 287940 306348 287946 306400
rect 288710 306348 288716 306400
rect 288768 306388 288774 306400
rect 289538 306388 289544 306400
rect 288768 306360 289544 306388
rect 288768 306348 288774 306360
rect 289538 306348 289544 306360
rect 289596 306348 289602 306400
rect 290182 306348 290188 306400
rect 290240 306388 290246 306400
rect 290826 306388 290832 306400
rect 290240 306360 290832 306388
rect 290240 306348 290246 306360
rect 290826 306348 290832 306360
rect 290884 306348 290890 306400
rect 292574 306348 292580 306400
rect 292632 306388 292638 306400
rect 293034 306388 293040 306400
rect 292632 306360 293040 306388
rect 292632 306348 292638 306360
rect 293034 306348 293040 306360
rect 293092 306348 293098 306400
rect 294046 306348 294052 306400
rect 294104 306388 294110 306400
rect 294322 306388 294328 306400
rect 294104 306360 294328 306388
rect 294104 306348 294110 306360
rect 294322 306348 294328 306360
rect 294380 306348 294386 306400
rect 295334 306348 295340 306400
rect 295392 306388 295398 306400
rect 295978 306388 295984 306400
rect 295392 306360 295984 306388
rect 295392 306348 295398 306360
rect 295978 306348 295984 306360
rect 296036 306348 296042 306400
rect 298094 306348 298100 306400
rect 298152 306388 298158 306400
rect 298554 306388 298560 306400
rect 298152 306360 298560 306388
rect 298152 306348 298158 306360
rect 298554 306348 298560 306360
rect 298612 306348 298618 306400
rect 301038 306348 301044 306400
rect 301096 306388 301102 306400
rect 301498 306388 301504 306400
rect 301096 306360 301504 306388
rect 301096 306348 301102 306360
rect 301498 306348 301504 306360
rect 301556 306348 301562 306400
rect 311894 306348 311900 306400
rect 311952 306388 311958 306400
rect 312170 306388 312176 306400
rect 311952 306360 312176 306388
rect 311952 306348 311958 306360
rect 312170 306348 312176 306360
rect 312228 306348 312234 306400
rect 313366 306348 313372 306400
rect 313424 306388 313430 306400
rect 314010 306388 314016 306400
rect 313424 306360 314016 306388
rect 313424 306348 313430 306360
rect 314010 306348 314016 306360
rect 314068 306348 314074 306400
rect 314654 306348 314660 306400
rect 314712 306388 314718 306400
rect 315114 306388 315120 306400
rect 314712 306360 315120 306388
rect 314712 306348 314718 306360
rect 315114 306348 315120 306360
rect 315172 306348 315178 306400
rect 317506 306348 317512 306400
rect 317564 306388 317570 306400
rect 318242 306388 318248 306400
rect 317564 306360 318248 306388
rect 317564 306348 317570 306360
rect 318242 306348 318248 306360
rect 318300 306348 318306 306400
rect 318886 306348 318892 306400
rect 318944 306388 318950 306400
rect 319530 306388 319536 306400
rect 318944 306360 319536 306388
rect 318944 306348 318950 306360
rect 319530 306348 319536 306360
rect 319588 306348 319594 306400
rect 320174 306348 320180 306400
rect 320232 306388 320238 306400
rect 321002 306388 321008 306400
rect 320232 306360 321008 306388
rect 320232 306348 320238 306360
rect 321002 306348 321008 306360
rect 321060 306348 321066 306400
rect 321554 306348 321560 306400
rect 321612 306388 321618 306400
rect 321922 306388 321928 306400
rect 321612 306360 321928 306388
rect 321612 306348 321618 306360
rect 321922 306348 321928 306360
rect 321980 306348 321986 306400
rect 326062 306348 326068 306400
rect 326120 306388 326126 306400
rect 326522 306388 326528 306400
rect 326120 306360 326528 306388
rect 326120 306348 326126 306360
rect 326522 306348 326528 306360
rect 326580 306348 326586 306400
rect 327166 306348 327172 306400
rect 327224 306388 327230 306400
rect 327810 306388 327816 306400
rect 327224 306360 327816 306388
rect 327224 306348 327230 306360
rect 327810 306348 327816 306360
rect 327868 306348 327874 306400
rect 328822 306348 328828 306400
rect 328880 306388 328886 306400
rect 329098 306388 329104 306400
rect 328880 306360 329104 306388
rect 328880 306348 328886 306360
rect 329098 306348 329104 306360
rect 329156 306348 329162 306400
rect 331490 306348 331496 306400
rect 331548 306388 331554 306400
rect 332410 306388 332416 306400
rect 331548 306360 332416 306388
rect 331548 306348 331554 306360
rect 332410 306348 332416 306360
rect 332468 306348 332474 306400
rect 341058 306348 341064 306400
rect 341116 306388 341122 306400
rect 341334 306388 341340 306400
rect 341116 306360 341340 306388
rect 341116 306348 341122 306360
rect 341334 306348 341340 306360
rect 341392 306348 341398 306400
rect 347958 306348 347964 306400
rect 348016 306348 348022 306400
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 228358 306320 228364 306332
rect 3384 306292 228364 306320
rect 3384 306280 3390 306292
rect 228358 306280 228364 306292
rect 228416 306280 228422 306332
rect 255406 306280 255412 306332
rect 255464 306320 255470 306332
rect 256418 306320 256424 306332
rect 255464 306292 256424 306320
rect 255464 306280 255470 306292
rect 256418 306280 256424 306292
rect 256476 306280 256482 306332
rect 259822 306280 259828 306332
rect 259880 306320 259886 306332
rect 260650 306320 260656 306332
rect 259880 306292 260656 306320
rect 259880 306280 259886 306292
rect 260650 306280 260656 306292
rect 260708 306280 260714 306332
rect 260926 306280 260932 306332
rect 260984 306320 260990 306332
rect 261570 306320 261576 306332
rect 260984 306292 261576 306320
rect 260984 306280 260990 306292
rect 261570 306280 261576 306292
rect 261628 306280 261634 306332
rect 262582 306280 262588 306332
rect 262640 306320 262646 306332
rect 262858 306320 262864 306332
rect 262640 306292 262864 306320
rect 262640 306280 262646 306292
rect 262858 306280 262864 306292
rect 262916 306280 262922 306332
rect 273346 306280 273352 306332
rect 273404 306320 273410 306332
rect 274082 306320 274088 306332
rect 273404 306292 274088 306320
rect 273404 306280 273410 306292
rect 274082 306280 274088 306292
rect 274140 306280 274146 306332
rect 274818 306280 274824 306332
rect 274876 306320 274882 306332
rect 275738 306320 275744 306332
rect 274876 306292 275744 306320
rect 274876 306280 274882 306292
rect 275738 306280 275744 306292
rect 275796 306280 275802 306332
rect 276106 306280 276112 306332
rect 276164 306320 276170 306332
rect 276658 306320 276664 306332
rect 276164 306292 276664 306320
rect 276164 306280 276170 306292
rect 276658 306280 276664 306292
rect 276716 306280 276722 306332
rect 277578 306280 277584 306332
rect 277636 306320 277642 306332
rect 278682 306320 278688 306332
rect 277636 306292 278688 306320
rect 277636 306280 277642 306292
rect 278682 306280 278688 306292
rect 278740 306280 278746 306332
rect 280338 306280 280344 306332
rect 280396 306320 280402 306332
rect 281074 306320 281080 306332
rect 280396 306292 281080 306320
rect 280396 306280 280402 306292
rect 281074 306280 281080 306292
rect 281132 306280 281138 306332
rect 281902 306280 281908 306332
rect 281960 306320 281966 306332
rect 282178 306320 282184 306332
rect 281960 306292 282184 306320
rect 281960 306280 281966 306292
rect 282178 306280 282184 306292
rect 282236 306280 282242 306332
rect 282270 306280 282276 306332
rect 282328 306320 282334 306332
rect 334802 306320 334808 306332
rect 282328 306292 334808 306320
rect 282328 306280 282334 306292
rect 334802 306280 334808 306292
rect 334860 306280 334866 306332
rect 254210 306212 254216 306264
rect 254268 306252 254274 306264
rect 254762 306252 254768 306264
rect 254268 306224 254768 306252
rect 254268 306212 254274 306224
rect 254762 306212 254768 306224
rect 254820 306212 254826 306264
rect 256786 306212 256792 306264
rect 256844 306252 256850 306264
rect 257522 306252 257528 306264
rect 256844 306224 257528 306252
rect 256844 306212 256850 306224
rect 257522 306212 257528 306224
rect 257580 306212 257586 306264
rect 258166 306212 258172 306264
rect 258224 306252 258230 306264
rect 259362 306252 259368 306264
rect 258224 306224 259368 306252
rect 258224 306212 258230 306224
rect 259362 306212 259368 306224
rect 259420 306212 259426 306264
rect 259638 306212 259644 306264
rect 259696 306252 259702 306264
rect 260006 306252 260012 306264
rect 259696 306224 260012 306252
rect 259696 306212 259702 306224
rect 260006 306212 260012 306224
rect 260064 306212 260070 306264
rect 260834 306212 260840 306264
rect 260892 306252 260898 306264
rect 261294 306252 261300 306264
rect 260892 306224 261300 306252
rect 260892 306212 260898 306224
rect 261294 306212 261300 306224
rect 261352 306212 261358 306264
rect 262490 306212 262496 306264
rect 262548 306252 262554 306264
rect 263410 306252 263416 306264
rect 262548 306224 263416 306252
rect 262548 306212 262554 306224
rect 263410 306212 263416 306224
rect 263468 306212 263474 306264
rect 271782 306212 271788 306264
rect 271840 306252 271846 306264
rect 329374 306252 329380 306264
rect 271840 306224 329380 306252
rect 271840 306212 271846 306224
rect 329374 306212 329380 306224
rect 329432 306212 329438 306264
rect 334158 306212 334164 306264
rect 334216 306252 334222 306264
rect 335170 306252 335176 306264
rect 334216 306224 335176 306252
rect 334216 306212 334222 306224
rect 335170 306212 335176 306224
rect 335228 306212 335234 306264
rect 335354 306212 335360 306264
rect 335412 306252 335418 306264
rect 335814 306252 335820 306264
rect 335412 306224 335820 306252
rect 335412 306212 335418 306224
rect 335814 306212 335820 306224
rect 335872 306212 335878 306264
rect 336918 306212 336924 306264
rect 336976 306252 336982 306264
rect 337562 306252 337568 306264
rect 336976 306224 337568 306252
rect 336976 306212 336982 306224
rect 337562 306212 337568 306224
rect 337620 306212 337626 306264
rect 338298 306212 338304 306264
rect 338356 306252 338362 306264
rect 339218 306252 339224 306264
rect 338356 306224 339224 306252
rect 338356 306212 338362 306224
rect 339218 306212 339224 306224
rect 339276 306212 339282 306264
rect 339678 306212 339684 306264
rect 339736 306252 339742 306264
rect 340506 306252 340512 306264
rect 339736 306224 340512 306252
rect 339736 306212 339742 306224
rect 340506 306212 340512 306224
rect 340564 306212 340570 306264
rect 256878 306144 256884 306196
rect 256936 306184 256942 306196
rect 257890 306184 257896 306196
rect 256936 306156 257896 306184
rect 256936 306144 256942 306156
rect 257890 306144 257896 306156
rect 257948 306144 257954 306196
rect 275002 306144 275008 306196
rect 275060 306184 275066 306196
rect 275554 306184 275560 306196
rect 275060 306156 275560 306184
rect 275060 306144 275066 306156
rect 275554 306144 275560 306156
rect 275612 306144 275618 306196
rect 276474 306144 276480 306196
rect 276532 306184 276538 306196
rect 277026 306184 277032 306196
rect 276532 306156 277032 306184
rect 276532 306144 276538 306156
rect 277026 306144 277032 306156
rect 277084 306144 277090 306196
rect 280522 306144 280528 306196
rect 280580 306184 280586 306196
rect 281442 306184 281448 306196
rect 280580 306156 281448 306184
rect 280580 306144 280586 306156
rect 281442 306144 281448 306156
rect 281500 306144 281506 306196
rect 281534 306144 281540 306196
rect 281592 306184 281598 306196
rect 281592 306156 332364 306184
rect 281592 306144 281598 306156
rect 255314 306076 255320 306128
rect 255372 306116 255378 306128
rect 255866 306116 255872 306128
rect 255372 306088 255872 306116
rect 255372 306076 255378 306088
rect 255866 306076 255872 306088
rect 255924 306076 255930 306128
rect 257154 306076 257160 306128
rect 257212 306116 257218 306128
rect 257706 306116 257712 306128
rect 257212 306088 257712 306116
rect 257212 306076 257218 306088
rect 257706 306076 257712 306088
rect 257764 306076 257770 306128
rect 259638 306076 259644 306128
rect 259696 306116 259702 306128
rect 260282 306116 260288 306128
rect 259696 306088 260288 306116
rect 259696 306076 259702 306088
rect 260282 306076 260288 306088
rect 260340 306076 260346 306128
rect 260834 306076 260840 306128
rect 260892 306116 260898 306128
rect 262122 306116 262128 306128
rect 260892 306088 262128 306116
rect 260892 306076 260898 306088
rect 262122 306076 262128 306088
rect 262180 306076 262186 306128
rect 271690 306076 271696 306128
rect 271748 306116 271754 306128
rect 332226 306116 332232 306128
rect 271748 306088 332232 306116
rect 271748 306076 271754 306088
rect 332226 306076 332232 306088
rect 332284 306076 332290 306128
rect 332336 306116 332364 306156
rect 335538 306116 335544 306128
rect 332336 306088 335544 306116
rect 335538 306076 335544 306088
rect 335596 306076 335602 306128
rect 273622 306008 273628 306060
rect 273680 306048 273686 306060
rect 274450 306048 274456 306060
rect 273680 306020 274456 306048
rect 273680 306008 273686 306020
rect 274450 306008 274456 306020
rect 274508 306008 274514 306060
rect 276290 306008 276296 306060
rect 276348 306048 276354 306060
rect 276842 306048 276848 306060
rect 276348 306020 276848 306048
rect 276348 306008 276354 306020
rect 276842 306008 276848 306020
rect 276900 306008 276906 306060
rect 277762 306008 277768 306060
rect 277820 306048 277826 306060
rect 278498 306048 278504 306060
rect 277820 306020 278504 306048
rect 277820 306008 277826 306020
rect 278498 306008 278504 306020
rect 278556 306008 278562 306060
rect 278590 306008 278596 306060
rect 278648 306048 278654 306060
rect 344554 306048 344560 306060
rect 278648 306020 344560 306048
rect 278648 306008 278654 306020
rect 344554 306008 344560 306020
rect 344612 306008 344618 306060
rect 255590 305940 255596 305992
rect 255648 305980 255654 305992
rect 256602 305980 256608 305992
rect 255648 305952 256608 305980
rect 255648 305940 255654 305952
rect 256602 305940 256608 305952
rect 256660 305940 256666 305992
rect 256970 305940 256976 305992
rect 257028 305980 257034 305992
rect 257338 305980 257344 305992
rect 257028 305952 257344 305980
rect 257028 305940 257034 305952
rect 257338 305940 257344 305952
rect 257396 305940 257402 305992
rect 275278 305940 275284 305992
rect 275336 305980 275342 305992
rect 345014 305980 345020 305992
rect 275336 305952 345020 305980
rect 275336 305940 275342 305952
rect 345014 305940 345020 305952
rect 345072 305940 345078 305992
rect 255682 305872 255688 305924
rect 255740 305912 255746 305924
rect 256234 305912 256240 305924
rect 255740 305884 256240 305912
rect 255740 305872 255746 305884
rect 256234 305872 256240 305884
rect 256292 305872 256298 305924
rect 272610 305872 272616 305924
rect 272668 305912 272674 305924
rect 345106 305912 345112 305924
rect 272668 305884 345112 305912
rect 272668 305872 272674 305884
rect 345106 305872 345112 305884
rect 345164 305872 345170 305924
rect 272518 305804 272524 305856
rect 272576 305844 272582 305856
rect 345198 305844 345204 305856
rect 272576 305816 345204 305844
rect 272576 305804 272582 305816
rect 345198 305804 345204 305816
rect 345256 305804 345262 305856
rect 88978 305736 88984 305788
rect 89036 305776 89042 305788
rect 253290 305776 253296 305788
rect 89036 305748 253296 305776
rect 89036 305736 89042 305748
rect 253290 305736 253296 305748
rect 253348 305736 253354 305788
rect 269850 305736 269856 305788
rect 269908 305776 269914 305788
rect 347314 305776 347320 305788
rect 269908 305748 347320 305776
rect 269908 305736 269914 305748
rect 347314 305736 347320 305748
rect 347372 305736 347378 305788
rect 71774 305668 71780 305720
rect 71832 305708 71838 305720
rect 251266 305708 251272 305720
rect 71832 305680 251272 305708
rect 71832 305668 71838 305680
rect 251266 305668 251272 305680
rect 251324 305668 251330 305720
rect 270034 305668 270040 305720
rect 270092 305708 270098 305720
rect 347774 305708 347780 305720
rect 270092 305680 347780 305708
rect 270092 305668 270098 305680
rect 347774 305668 347780 305680
rect 347832 305668 347838 305720
rect 35158 305600 35164 305652
rect 35216 305640 35222 305652
rect 244458 305640 244464 305652
rect 35216 305612 244464 305640
rect 35216 305600 35222 305612
rect 244458 305600 244464 305612
rect 244516 305600 244522 305652
rect 266998 305600 267004 305652
rect 267056 305640 267062 305652
rect 347866 305640 347872 305652
rect 267056 305612 347872 305640
rect 267056 305600 267062 305612
rect 347866 305600 347872 305612
rect 347924 305600 347930 305652
rect 257338 305532 257344 305584
rect 257396 305572 257402 305584
rect 257982 305572 257988 305584
rect 257396 305544 257988 305572
rect 257396 305532 257402 305544
rect 257982 305532 257988 305544
rect 258040 305532 258046 305584
rect 275370 305532 275376 305584
rect 275428 305572 275434 305584
rect 278590 305572 278596 305584
rect 275428 305544 278596 305572
rect 275428 305532 275434 305544
rect 278590 305532 278596 305544
rect 278648 305532 278654 305584
rect 279418 305532 279424 305584
rect 279476 305572 279482 305584
rect 279878 305572 279884 305584
rect 279476 305544 279884 305572
rect 279476 305532 279482 305544
rect 279878 305532 279884 305544
rect 279936 305532 279942 305584
rect 281442 305532 281448 305584
rect 281500 305572 281506 305584
rect 281500 305544 332364 305572
rect 281500 305532 281506 305544
rect 274542 305464 274548 305516
rect 274600 305504 274606 305516
rect 281534 305504 281540 305516
rect 274600 305476 281540 305504
rect 274600 305464 274606 305476
rect 281534 305464 281540 305476
rect 281592 305464 281598 305516
rect 284570 305464 284576 305516
rect 284628 305504 284634 305516
rect 284938 305504 284944 305516
rect 284628 305476 284944 305504
rect 284628 305464 284634 305476
rect 284938 305464 284944 305476
rect 284996 305464 285002 305516
rect 285858 305464 285864 305516
rect 285916 305504 285922 305516
rect 286962 305504 286968 305516
rect 285916 305476 286968 305504
rect 285916 305464 285922 305476
rect 286962 305464 286968 305476
rect 287020 305464 287026 305516
rect 287146 305464 287152 305516
rect 287204 305504 287210 305516
rect 287514 305504 287520 305516
rect 287204 305476 287520 305504
rect 287204 305464 287210 305476
rect 287514 305464 287520 305476
rect 287572 305464 287578 305516
rect 288434 305464 288440 305516
rect 288492 305504 288498 305516
rect 288894 305504 288900 305516
rect 288492 305476 288900 305504
rect 288492 305464 288498 305476
rect 288894 305464 288900 305476
rect 288952 305464 288958 305516
rect 290090 305464 290096 305516
rect 290148 305504 290154 305516
rect 290642 305504 290648 305516
rect 290148 305476 290648 305504
rect 290148 305464 290154 305476
rect 290642 305464 290648 305476
rect 290700 305464 290706 305516
rect 291378 305464 291384 305516
rect 291436 305504 291442 305516
rect 291746 305504 291752 305516
rect 291436 305476 291752 305504
rect 291436 305464 291442 305476
rect 291746 305464 291752 305476
rect 291804 305464 291810 305516
rect 292390 305464 292396 305516
rect 292448 305504 292454 305516
rect 292448 305476 332272 305504
rect 292448 305464 292454 305476
rect 274358 305396 274364 305448
rect 274416 305436 274422 305448
rect 282270 305436 282276 305448
rect 274416 305408 282276 305436
rect 274416 305396 274422 305408
rect 282270 305396 282276 305408
rect 282328 305396 282334 305448
rect 288618 305396 288624 305448
rect 288676 305436 288682 305448
rect 289722 305436 289728 305448
rect 288676 305408 289728 305436
rect 288676 305396 288682 305408
rect 289722 305396 289728 305408
rect 289780 305396 289786 305448
rect 289906 305396 289912 305448
rect 289964 305436 289970 305448
rect 290458 305436 290464 305448
rect 289964 305408 290464 305436
rect 289964 305396 289970 305408
rect 290458 305396 290464 305408
rect 290516 305396 290522 305448
rect 291562 305396 291568 305448
rect 291620 305436 291626 305448
rect 292114 305436 292120 305448
rect 291620 305408 292120 305436
rect 291620 305396 291626 305408
rect 292114 305396 292120 305408
rect 292172 305396 292178 305448
rect 294046 305396 294052 305448
rect 294104 305436 294110 305448
rect 295058 305436 295064 305448
rect 294104 305408 295064 305436
rect 294104 305396 294110 305408
rect 295058 305396 295064 305408
rect 295116 305396 295122 305448
rect 295518 305396 295524 305448
rect 295576 305436 295582 305448
rect 296162 305436 296168 305448
rect 295576 305408 296168 305436
rect 295576 305396 295582 305408
rect 296162 305396 296168 305408
rect 296220 305396 296226 305448
rect 296990 305396 296996 305448
rect 297048 305436 297054 305448
rect 297634 305436 297640 305448
rect 297048 305408 297640 305436
rect 297048 305396 297054 305408
rect 297634 305396 297640 305408
rect 297692 305396 297698 305448
rect 298370 305396 298376 305448
rect 298428 305436 298434 305448
rect 299290 305436 299296 305448
rect 298428 305408 299296 305436
rect 298428 305396 298434 305408
rect 299290 305396 299296 305408
rect 299348 305396 299354 305448
rect 299658 305396 299664 305448
rect 299716 305436 299722 305448
rect 300026 305436 300032 305448
rect 299716 305408 300032 305436
rect 299716 305396 299722 305408
rect 300026 305396 300032 305408
rect 300084 305396 300090 305448
rect 301222 305396 301228 305448
rect 301280 305436 301286 305448
rect 301866 305436 301872 305448
rect 301280 305408 301872 305436
rect 301280 305396 301286 305408
rect 301866 305396 301872 305408
rect 301924 305396 301930 305448
rect 332042 305436 332048 305448
rect 302206 305408 332048 305436
rect 278038 305328 278044 305380
rect 278096 305368 278102 305380
rect 278222 305368 278228 305380
rect 278096 305340 278228 305368
rect 278096 305328 278102 305340
rect 278222 305328 278228 305340
rect 278280 305328 278286 305380
rect 287146 305328 287152 305380
rect 287204 305368 287210 305380
rect 288066 305368 288072 305380
rect 287204 305340 288072 305368
rect 287204 305328 287210 305340
rect 288066 305328 288072 305340
rect 288124 305328 288130 305380
rect 288434 305328 288440 305380
rect 288492 305368 288498 305380
rect 289170 305368 289176 305380
rect 288492 305340 289176 305368
rect 288492 305328 288498 305340
rect 289170 305328 289176 305340
rect 289228 305328 289234 305380
rect 291286 305328 291292 305380
rect 291344 305368 291350 305380
rect 292298 305368 292304 305380
rect 291344 305340 292304 305368
rect 291344 305328 291350 305340
rect 292298 305328 292304 305340
rect 292356 305328 292362 305380
rect 299566 305328 299572 305380
rect 299624 305368 299630 305380
rect 300578 305368 300584 305380
rect 299624 305340 300584 305368
rect 299624 305328 299630 305340
rect 300578 305328 300584 305340
rect 300636 305328 300642 305380
rect 301130 305328 301136 305380
rect 301188 305368 301194 305380
rect 301682 305368 301688 305380
rect 301188 305340 301688 305368
rect 301188 305328 301194 305340
rect 301682 305328 301688 305340
rect 301740 305328 301746 305380
rect 277946 305260 277952 305312
rect 278004 305300 278010 305312
rect 278314 305300 278320 305312
rect 278004 305272 278320 305300
rect 278004 305260 278010 305272
rect 278314 305260 278320 305272
rect 278372 305260 278378 305312
rect 299474 305260 299480 305312
rect 299532 305300 299538 305312
rect 300394 305300 300400 305312
rect 299532 305272 300400 305300
rect 299532 305260 299538 305272
rect 300394 305260 300400 305272
rect 300452 305260 300458 305312
rect 298278 305192 298284 305244
rect 298336 305232 298342 305244
rect 298738 305232 298744 305244
rect 298336 305204 298744 305232
rect 298336 305192 298342 305204
rect 298738 305192 298744 305204
rect 298796 305192 298802 305244
rect 302206 305232 302234 305408
rect 332042 305396 332048 305408
rect 332100 305396 332106 305448
rect 313642 305328 313648 305380
rect 313700 305368 313706 305380
rect 313826 305368 313832 305380
rect 313700 305340 313832 305368
rect 313700 305328 313706 305340
rect 313826 305328 313832 305340
rect 313884 305328 313890 305380
rect 316034 305328 316040 305380
rect 316092 305368 316098 305380
rect 316402 305368 316408 305380
rect 316092 305340 316408 305368
rect 316092 305328 316098 305340
rect 316402 305328 316408 305340
rect 316460 305328 316466 305380
rect 317782 305328 317788 305380
rect 317840 305368 317846 305380
rect 318610 305368 318616 305380
rect 317840 305340 318616 305368
rect 317840 305328 317846 305340
rect 318610 305328 318616 305340
rect 318668 305328 318674 305380
rect 318978 305328 318984 305380
rect 319036 305368 319042 305380
rect 319254 305368 319260 305380
rect 319036 305340 319260 305368
rect 319036 305328 319042 305340
rect 319254 305328 319260 305340
rect 319312 305328 319318 305380
rect 320542 305328 320548 305380
rect 320600 305368 320606 305380
rect 321370 305368 321376 305380
rect 320600 305340 321376 305368
rect 320600 305328 320606 305340
rect 321370 305328 321376 305340
rect 321428 305328 321434 305380
rect 321830 305328 321836 305380
rect 321888 305368 321894 305380
rect 322290 305368 322296 305380
rect 321888 305340 322296 305368
rect 321888 305328 321894 305340
rect 322290 305328 322296 305340
rect 322348 305328 322354 305380
rect 323302 305328 323308 305380
rect 323360 305368 323366 305380
rect 324130 305368 324136 305380
rect 323360 305340 324136 305368
rect 323360 305328 323366 305340
rect 324130 305328 324136 305340
rect 324188 305328 324194 305380
rect 324314 305328 324320 305380
rect 324372 305368 324378 305380
rect 324590 305368 324596 305380
rect 324372 305340 324596 305368
rect 324372 305328 324378 305340
rect 324590 305328 324596 305340
rect 324648 305328 324654 305380
rect 324866 305328 324872 305380
rect 324924 305368 324930 305380
rect 325602 305368 325608 305380
rect 324924 305340 325608 305368
rect 324924 305328 324930 305340
rect 325602 305328 325608 305340
rect 325660 305328 325666 305380
rect 326154 305328 326160 305380
rect 326212 305368 326218 305380
rect 326706 305368 326712 305380
rect 326212 305340 326712 305368
rect 326212 305328 326218 305340
rect 326706 305328 326712 305340
rect 326764 305328 326770 305380
rect 327074 305328 327080 305380
rect 327132 305368 327138 305380
rect 327626 305368 327632 305380
rect 327132 305340 327632 305368
rect 327132 305328 327138 305340
rect 327626 305328 327632 305340
rect 327684 305328 327690 305380
rect 328730 305328 328736 305380
rect 328788 305368 328794 305380
rect 329650 305368 329656 305380
rect 328788 305340 329656 305368
rect 328788 305328 328794 305340
rect 329650 305328 329656 305340
rect 329708 305328 329714 305380
rect 332244 305368 332272 305476
rect 332336 305436 332364 305544
rect 332410 305532 332416 305584
rect 332468 305572 332474 305584
rect 337194 305572 337200 305584
rect 332468 305544 337200 305572
rect 332468 305532 332474 305544
rect 337194 305532 337200 305544
rect 337252 305532 337258 305584
rect 336274 305436 336280 305448
rect 332336 305408 336280 305436
rect 336274 305396 336280 305408
rect 336332 305396 336338 305448
rect 333882 305368 333888 305380
rect 332244 305340 333888 305368
rect 333882 305328 333888 305340
rect 333940 305328 333946 305380
rect 316310 305260 316316 305312
rect 316368 305300 316374 305312
rect 317138 305300 317144 305312
rect 316368 305272 317144 305300
rect 316368 305260 316374 305272
rect 317138 305260 317144 305272
rect 317196 305260 317202 305312
rect 318794 305260 318800 305312
rect 318852 305300 318858 305312
rect 319162 305300 319168 305312
rect 318852 305272 319168 305300
rect 318852 305260 318858 305272
rect 319162 305260 319168 305272
rect 319220 305260 319226 305312
rect 320358 305260 320364 305312
rect 320416 305300 320422 305312
rect 321186 305300 321192 305312
rect 320416 305272 321192 305300
rect 320416 305260 320422 305272
rect 321186 305260 321192 305272
rect 321244 305260 321250 305312
rect 321646 305260 321652 305312
rect 321704 305300 321710 305312
rect 322474 305300 322480 305312
rect 321704 305272 322480 305300
rect 321704 305260 321710 305272
rect 322474 305260 322480 305272
rect 322532 305260 322538 305312
rect 322934 305260 322940 305312
rect 322992 305300 322998 305312
rect 323486 305300 323492 305312
rect 322992 305272 323492 305300
rect 322992 305260 322998 305272
rect 323486 305260 323492 305272
rect 323544 305260 323550 305312
rect 325786 305260 325792 305312
rect 325844 305300 325850 305312
rect 326890 305300 326896 305312
rect 325844 305272 326896 305300
rect 325844 305260 325850 305272
rect 326890 305260 326896 305272
rect 326948 305260 326954 305312
rect 327258 305260 327264 305312
rect 327316 305300 327322 305312
rect 328362 305300 328368 305312
rect 327316 305272 328368 305300
rect 327316 305260 327322 305272
rect 328362 305260 328368 305272
rect 328420 305260 328426 305312
rect 328546 305260 328552 305312
rect 328604 305300 328610 305312
rect 329282 305300 329288 305312
rect 328604 305272 329288 305300
rect 328604 305260 328610 305272
rect 329282 305260 329288 305272
rect 329340 305260 329346 305312
rect 298848 305204 302234 305232
rect 296530 305124 296536 305176
rect 296588 305164 296594 305176
rect 298848 305164 298876 305204
rect 316402 305192 316408 305244
rect 316460 305232 316466 305244
rect 317322 305232 317328 305244
rect 316460 305204 317328 305232
rect 316460 305192 316466 305204
rect 317322 305192 317328 305204
rect 317380 305192 317386 305244
rect 318978 305192 318984 305244
rect 319036 305232 319042 305244
rect 319898 305232 319904 305244
rect 319036 305204 319904 305232
rect 319036 305192 319042 305204
rect 319898 305192 319904 305204
rect 319956 305192 319962 305244
rect 321738 305192 321744 305244
rect 321796 305232 321802 305244
rect 322842 305232 322848 305244
rect 321796 305204 322848 305232
rect 321796 305192 321802 305204
rect 322842 305192 322848 305204
rect 322900 305192 322906 305244
rect 323210 305192 323216 305244
rect 323268 305232 323274 305244
rect 323946 305232 323952 305244
rect 323268 305204 323952 305232
rect 323268 305192 323274 305204
rect 323946 305192 323952 305204
rect 324004 305192 324010 305244
rect 324590 305192 324596 305244
rect 324648 305232 324654 305244
rect 325418 305232 325424 305244
rect 324648 305204 325424 305232
rect 324648 305192 324654 305204
rect 325418 305192 325424 305204
rect 325476 305192 325482 305244
rect 327074 305192 327080 305244
rect 327132 305232 327138 305244
rect 328178 305232 328184 305244
rect 327132 305204 328184 305232
rect 327132 305192 327138 305204
rect 328178 305192 328184 305204
rect 328236 305192 328242 305244
rect 296588 305136 298876 305164
rect 296588 305124 296594 305136
rect 299934 305124 299940 305176
rect 299992 305164 299998 305176
rect 300762 305164 300768 305176
rect 299992 305136 300768 305164
rect 299992 305124 299998 305136
rect 300762 305124 300768 305136
rect 300820 305124 300826 305176
rect 318794 305124 318800 305176
rect 318852 305164 318858 305176
rect 320082 305164 320088 305176
rect 318852 305136 320088 305164
rect 318852 305124 318858 305136
rect 320082 305124 320088 305136
rect 320140 305124 320146 305176
rect 322106 305124 322112 305176
rect 322164 305164 322170 305176
rect 322658 305164 322664 305176
rect 322164 305136 322664 305164
rect 322164 305124 322170 305136
rect 322658 305124 322664 305136
rect 322716 305124 322722 305176
rect 322934 305124 322940 305176
rect 322992 305164 322998 305176
rect 323762 305164 323768 305176
rect 322992 305136 323768 305164
rect 322992 305124 322998 305136
rect 323762 305124 323768 305136
rect 323820 305124 323826 305176
rect 282914 305056 282920 305108
rect 282972 305096 282978 305108
rect 284018 305096 284024 305108
rect 282972 305068 284024 305096
rect 282972 305056 282978 305068
rect 284018 305056 284024 305068
rect 284076 305056 284082 305108
rect 294138 305056 294144 305108
rect 294196 305096 294202 305108
rect 294506 305096 294512 305108
rect 294196 305068 294512 305096
rect 294196 305056 294202 305068
rect 294506 305056 294512 305068
rect 294564 305056 294570 305108
rect 296806 304920 296812 304972
rect 296864 304960 296870 304972
rect 297450 304960 297456 304972
rect 296864 304932 297456 304960
rect 296864 304920 296870 304932
rect 297450 304920 297456 304932
rect 297508 304920 297514 304972
rect 278866 304648 278872 304700
rect 278924 304688 278930 304700
rect 279970 304688 279976 304700
rect 278924 304660 279976 304688
rect 278924 304648 278930 304660
rect 279970 304648 279976 304660
rect 280028 304648 280034 304700
rect 313550 304580 313556 304632
rect 313608 304620 313614 304632
rect 314194 304620 314200 304632
rect 313608 304592 314200 304620
rect 313608 304580 313614 304592
rect 314194 304580 314200 304592
rect 314252 304580 314258 304632
rect 313458 304512 313464 304564
rect 313516 304552 313522 304564
rect 314378 304552 314384 304564
rect 313516 304524 314384 304552
rect 313516 304512 313522 304524
rect 314378 304512 314384 304524
rect 314436 304512 314442 304564
rect 91094 304376 91100 304428
rect 91152 304416 91158 304428
rect 253934 304416 253940 304428
rect 91152 304388 253940 304416
rect 91152 304376 91158 304388
rect 253934 304376 253940 304388
rect 253992 304376 253998 304428
rect 317414 304376 317420 304428
rect 317472 304416 317478 304428
rect 318426 304416 318432 304428
rect 317472 304388 318432 304416
rect 317472 304376 317478 304388
rect 318426 304376 318432 304388
rect 318484 304376 318490 304428
rect 18598 304308 18604 304360
rect 18656 304348 18662 304360
rect 241606 304348 241612 304360
rect 18656 304320 241612 304348
rect 18656 304308 18662 304320
rect 241606 304308 241612 304320
rect 241664 304308 241670 304360
rect 254394 304308 254400 304360
rect 254452 304348 254458 304360
rect 254578 304348 254584 304360
rect 254452 304320 254584 304348
rect 254452 304308 254458 304320
rect 254578 304308 254584 304320
rect 254636 304308 254642 304360
rect 315850 304308 315856 304360
rect 315908 304348 315914 304360
rect 485038 304348 485044 304360
rect 315908 304320 485044 304348
rect 315908 304308 315914 304320
rect 485038 304308 485044 304320
rect 485096 304308 485102 304360
rect 13078 304240 13084 304292
rect 13136 304280 13142 304292
rect 240226 304280 240232 304292
rect 13136 304252 240232 304280
rect 13136 304240 13142 304252
rect 240226 304240 240232 304252
rect 240284 304240 240290 304292
rect 254118 304240 254124 304292
rect 254176 304280 254182 304292
rect 255130 304280 255136 304292
rect 254176 304252 255136 304280
rect 254176 304240 254182 304252
rect 255130 304240 255136 304252
rect 255188 304240 255194 304292
rect 292482 304240 292488 304292
rect 292540 304280 292546 304292
rect 292942 304280 292948 304292
rect 292540 304252 292948 304280
rect 292540 304240 292546 304252
rect 292942 304240 292948 304252
rect 293000 304240 293006 304292
rect 319346 304240 319352 304292
rect 319404 304280 319410 304292
rect 507854 304280 507860 304292
rect 319404 304252 507860 304280
rect 319404 304240 319410 304252
rect 507854 304240 507860 304252
rect 507912 304240 507918 304292
rect 335630 303832 335636 303884
rect 335688 303872 335694 303884
rect 336642 303872 336648 303884
rect 335688 303844 336648 303872
rect 335688 303832 335694 303844
rect 336642 303832 336648 303844
rect 336700 303832 336706 303884
rect 312170 303764 312176 303816
rect 312228 303804 312234 303816
rect 312538 303804 312544 303816
rect 312228 303776 312544 303804
rect 312228 303764 312234 303776
rect 312538 303764 312544 303776
rect 312596 303764 312602 303816
rect 311986 303696 311992 303748
rect 312044 303736 312050 303748
rect 312722 303736 312728 303748
rect 312044 303708 312728 303736
rect 312044 303696 312050 303708
rect 312722 303696 312728 303708
rect 312780 303696 312786 303748
rect 312078 303628 312084 303680
rect 312136 303668 312142 303680
rect 313090 303668 313096 303680
rect 312136 303640 313096 303668
rect 312136 303628 312142 303640
rect 313090 303628 313096 303640
rect 313148 303628 313154 303680
rect 282638 303560 282644 303612
rect 282696 303600 282702 303612
rect 330754 303600 330760 303612
rect 282696 303572 330760 303600
rect 282696 303560 282702 303572
rect 330754 303560 330760 303572
rect 330812 303560 330818 303612
rect 271598 303492 271604 303544
rect 271656 303532 271662 303544
rect 337746 303532 337752 303544
rect 271656 303504 337752 303532
rect 271656 303492 271662 303504
rect 337746 303492 337752 303504
rect 337804 303492 337810 303544
rect 261662 303424 261668 303476
rect 261720 303464 261726 303476
rect 334986 303464 334992 303476
rect 261720 303436 334992 303464
rect 261720 303424 261726 303436
rect 334986 303424 334992 303436
rect 335044 303424 335050 303476
rect 258902 303356 258908 303408
rect 258960 303396 258966 303408
rect 335538 303396 335544 303408
rect 258960 303368 335544 303396
rect 258960 303356 258966 303368
rect 335538 303356 335544 303368
rect 335596 303356 335602 303408
rect 258810 303288 258816 303340
rect 258868 303328 258874 303340
rect 336458 303328 336464 303340
rect 258868 303300 336464 303328
rect 258868 303288 258874 303300
rect 336458 303288 336464 303300
rect 336516 303288 336522 303340
rect 338390 303288 338396 303340
rect 338448 303328 338454 303340
rect 338666 303328 338672 303340
rect 338448 303300 338672 303328
rect 338448 303288 338454 303300
rect 338666 303288 338672 303300
rect 338724 303288 338730 303340
rect 258718 303220 258724 303272
rect 258776 303260 258782 303272
rect 337286 303260 337292 303272
rect 258776 303232 337292 303260
rect 258776 303220 258782 303232
rect 337286 303220 337292 303232
rect 337344 303220 337350 303272
rect 256142 303152 256148 303204
rect 256200 303192 256206 303204
rect 337930 303192 337936 303204
rect 256200 303164 337936 303192
rect 256200 303152 256206 303164
rect 337930 303152 337936 303164
rect 337988 303152 337994 303204
rect 267182 303084 267188 303136
rect 267240 303124 267246 303136
rect 348970 303124 348976 303136
rect 267240 303096 348976 303124
rect 267240 303084 267246 303096
rect 348970 303084 348976 303096
rect 349028 303084 349034 303136
rect 82814 303016 82820 303068
rect 82872 303056 82878 303068
rect 252646 303056 252652 303068
rect 82872 303028 252652 303056
rect 82872 303016 82878 303028
rect 252646 303016 252652 303028
rect 252704 303016 252710 303068
rect 256234 303016 256240 303068
rect 256292 303056 256298 303068
rect 338574 303056 338580 303068
rect 256292 303028 338580 303056
rect 256292 303016 256298 303028
rect 338574 303016 338580 303028
rect 338632 303016 338638 303068
rect 27614 302948 27620 303000
rect 27672 302988 27678 303000
rect 244642 302988 244648 303000
rect 27672 302960 244648 302988
rect 27672 302948 27678 302960
rect 244642 302948 244648 302960
rect 244700 302948 244706 303000
rect 264330 302948 264336 303000
rect 264388 302988 264394 303000
rect 349246 302988 349252 303000
rect 264388 302960 349252 302988
rect 264388 302948 264394 302960
rect 349246 302948 349252 302960
rect 349304 302948 349310 303000
rect 17218 302880 17224 302932
rect 17276 302920 17282 302932
rect 241146 302920 241152 302932
rect 17276 302892 241152 302920
rect 17276 302880 17282 302892
rect 241146 302880 241152 302892
rect 241204 302880 241210 302932
rect 261570 302880 261576 302932
rect 261628 302920 261634 302932
rect 350074 302920 350080 302932
rect 261628 302892 350080 302920
rect 261628 302880 261634 302892
rect 350074 302880 350080 302892
rect 350132 302880 350138 302932
rect 286686 302812 286692 302864
rect 286744 302852 286750 302864
rect 332594 302852 332600 302864
rect 286744 302824 332600 302852
rect 286744 302812 286750 302824
rect 332594 302812 332600 302824
rect 332652 302812 332658 302864
rect 283098 302744 283104 302796
rect 283156 302784 283162 302796
rect 283650 302784 283656 302796
rect 283156 302756 283656 302784
rect 283156 302744 283162 302756
rect 283650 302744 283656 302756
rect 283708 302744 283714 302796
rect 285490 302744 285496 302796
rect 285548 302784 285554 302796
rect 331674 302784 331680 302796
rect 285548 302756 331680 302784
rect 285548 302744 285554 302756
rect 331674 302744 331680 302756
rect 331732 302744 331738 302796
rect 293678 302676 293684 302728
rect 293736 302716 293742 302728
rect 331398 302716 331404 302728
rect 293736 302688 331404 302716
rect 293736 302676 293742 302688
rect 331398 302676 331404 302688
rect 331456 302676 331462 302728
rect 338114 302336 338120 302388
rect 338172 302376 338178 302388
rect 338574 302376 338580 302388
rect 338172 302348 338580 302376
rect 338172 302336 338178 302348
rect 338574 302336 338580 302348
rect 338632 302336 338638 302388
rect 294414 302200 294420 302252
rect 294472 302240 294478 302252
rect 294598 302240 294604 302252
rect 294472 302212 294604 302240
rect 294472 302200 294478 302212
rect 294598 302200 294604 302212
rect 294656 302200 294662 302252
rect 308490 301520 308496 301572
rect 308548 301560 308554 301572
rect 440234 301560 440240 301572
rect 308548 301532 440240 301560
rect 308548 301520 308554 301532
rect 440234 301520 440240 301532
rect 440292 301520 440298 301572
rect 39390 301452 39396 301504
rect 39448 301492 39454 301504
rect 245746 301492 245752 301504
rect 39448 301464 245752 301492
rect 39448 301452 39454 301464
rect 245746 301452 245752 301464
rect 245804 301452 245810 301504
rect 317874 301452 317880 301504
rect 317932 301492 317938 301504
rect 500218 301492 500224 301504
rect 317932 301464 500224 301492
rect 317932 301452 317938 301464
rect 500218 301452 500224 301464
rect 500276 301452 500282 301504
rect 289538 300704 289544 300756
rect 289596 300744 289602 300756
rect 334710 300744 334716 300756
rect 289596 300716 334716 300744
rect 289596 300704 289602 300716
rect 334710 300704 334716 300716
rect 334768 300704 334774 300756
rect 288066 300636 288072 300688
rect 288124 300676 288130 300688
rect 333514 300676 333520 300688
rect 288124 300648 333520 300676
rect 288124 300636 288130 300648
rect 333514 300636 333520 300648
rect 333572 300636 333578 300688
rect 286870 300568 286876 300620
rect 286928 300608 286934 300620
rect 333146 300608 333152 300620
rect 286928 300580 333152 300608
rect 286928 300568 286934 300580
rect 333146 300568 333152 300580
rect 333204 300568 333210 300620
rect 285398 300500 285404 300552
rect 285456 300540 285462 300552
rect 331490 300540 331496 300552
rect 285456 300512 331496 300540
rect 285456 300500 285462 300512
rect 331490 300500 331496 300512
rect 331548 300500 331554 300552
rect 284110 300432 284116 300484
rect 284168 300472 284174 300484
rect 341610 300472 341616 300484
rect 284168 300444 341616 300472
rect 284168 300432 284174 300444
rect 341610 300432 341616 300444
rect 341668 300432 341674 300484
rect 279970 300364 279976 300416
rect 280028 300404 280034 300416
rect 338850 300404 338856 300416
rect 280028 300376 338856 300404
rect 280028 300364 280034 300376
rect 338850 300364 338856 300376
rect 338908 300364 338914 300416
rect 277118 300296 277124 300348
rect 277176 300336 277182 300348
rect 339678 300336 339684 300348
rect 277176 300308 339684 300336
rect 277176 300296 277182 300308
rect 339678 300296 339684 300308
rect 339736 300296 339742 300348
rect 310146 300228 310152 300280
rect 310204 300268 310210 300280
rect 449894 300268 449900 300280
rect 310204 300240 449900 300268
rect 310204 300228 310210 300240
rect 449894 300228 449900 300240
rect 449952 300228 449958 300280
rect 71038 300160 71044 300212
rect 71096 300200 71102 300212
rect 249886 300200 249892 300212
rect 71096 300172 249892 300200
rect 71096 300160 71102 300172
rect 249886 300160 249892 300172
rect 249944 300160 249950 300212
rect 317782 300160 317788 300212
rect 317840 300200 317846 300212
rect 502978 300200 502984 300212
rect 317840 300172 502984 300200
rect 317840 300160 317846 300172
rect 502978 300160 502984 300172
rect 503036 300160 503042 300212
rect 21358 300092 21364 300144
rect 21416 300132 21422 300144
rect 242618 300132 242624 300144
rect 21416 300104 242624 300132
rect 21416 300092 21422 300104
rect 242618 300092 242624 300104
rect 242676 300092 242682 300144
rect 327626 300092 327632 300144
rect 327684 300132 327690 300144
rect 554038 300132 554044 300144
rect 327684 300104 554044 300132
rect 327684 300092 327690 300104
rect 554038 300092 554044 300104
rect 554096 300092 554102 300144
rect 70394 298868 70400 298920
rect 70452 298908 70458 298920
rect 251082 298908 251088 298920
rect 70452 298880 251088 298908
rect 70452 298868 70458 298880
rect 251082 298868 251088 298880
rect 251140 298868 251146 298920
rect 53834 298800 53840 298852
rect 53892 298840 53898 298852
rect 248506 298840 248512 298852
rect 53892 298812 248512 298840
rect 53892 298800 53898 298812
rect 248506 298800 248512 298812
rect 248564 298800 248570 298852
rect 312354 298800 312360 298852
rect 312412 298840 312418 298852
rect 462958 298840 462964 298852
rect 312412 298812 462964 298840
rect 312412 298800 312418 298812
rect 462958 298800 462964 298812
rect 463016 298800 463022 298852
rect 22738 298732 22744 298784
rect 22796 298772 22802 298784
rect 243170 298772 243176 298784
rect 22796 298744 243176 298772
rect 22796 298732 22802 298744
rect 243170 298732 243176 298744
rect 243228 298732 243234 298784
rect 319346 298732 319352 298784
rect 319404 298772 319410 298784
rect 511994 298772 512000 298784
rect 319404 298744 512000 298772
rect 319404 298732 319410 298744
rect 511994 298732 512000 298744
rect 512052 298732 512058 298784
rect 238294 297576 238300 297628
rect 238352 297616 238358 297628
rect 342898 297616 342904 297628
rect 238352 297588 342904 297616
rect 238352 297576 238358 297588
rect 342898 297576 342904 297588
rect 342956 297576 342962 297628
rect 92474 297508 92480 297560
rect 92532 297548 92538 297560
rect 254486 297548 254492 297560
rect 92532 297520 254492 297548
rect 92532 297508 92538 297520
rect 254486 297508 254492 297520
rect 254544 297508 254550 297560
rect 57974 297440 57980 297492
rect 58032 297480 58038 297492
rect 248782 297480 248788 297492
rect 58032 297452 248788 297480
rect 58032 297440 58038 297452
rect 248782 297440 248788 297452
rect 248840 297440 248846 297492
rect 35894 297372 35900 297424
rect 35952 297412 35958 297424
rect 246206 297412 246212 297424
rect 35952 297384 246212 297412
rect 35952 297372 35958 297384
rect 246206 297372 246212 297384
rect 246264 297372 246270 297424
rect 320634 297372 320640 297424
rect 320692 297412 320698 297424
rect 516778 297412 516784 297424
rect 320692 297384 516784 297412
rect 320692 297372 320698 297384
rect 516778 297372 516784 297384
rect 516836 297372 516842 297424
rect 80054 296012 80060 296064
rect 80112 296052 80118 296064
rect 253106 296052 253112 296064
rect 80112 296024 253112 296052
rect 80112 296012 80118 296024
rect 253106 296012 253112 296024
rect 253164 296012 253170 296064
rect 320542 296012 320548 296064
rect 320600 296052 320606 296064
rect 520918 296052 520924 296064
rect 320600 296024 520924 296052
rect 320600 296012 320606 296024
rect 520918 296012 520924 296024
rect 520976 296012 520982 296064
rect 60734 295944 60740 295996
rect 60792 295984 60798 295996
rect 248414 295984 248420 295996
rect 60792 295956 248420 295984
rect 60792 295944 60798 295956
rect 248414 295944 248420 295956
rect 248472 295944 248478 295996
rect 329006 295944 329012 295996
rect 329064 295984 329070 295996
rect 566458 295984 566464 295996
rect 329064 295956 566464 295984
rect 329064 295944 329070 295956
rect 566458 295944 566464 295956
rect 566516 295944 566522 295996
rect 310974 294788 310980 294840
rect 311032 294828 311038 294840
rect 453298 294828 453304 294840
rect 311032 294800 453304 294828
rect 311032 294788 311038 294800
rect 453298 294788 453304 294800
rect 453356 294788 453362 294840
rect 319254 294720 319260 294772
rect 319312 294760 319318 294772
rect 504358 294760 504364 294772
rect 319312 294732 504364 294760
rect 319312 294720 319318 294732
rect 504358 294720 504364 294732
rect 504416 294720 504422 294772
rect 69014 294652 69020 294704
rect 69072 294692 69078 294704
rect 250162 294692 250168 294704
rect 69072 294664 250168 294692
rect 69072 294652 69078 294664
rect 250162 294652 250168 294664
rect 250220 294652 250226 294704
rect 323486 294652 323492 294704
rect 323544 294692 323550 294704
rect 527818 294692 527824 294704
rect 323544 294664 527824 294692
rect 323544 294652 323550 294664
rect 527818 294652 527824 294664
rect 527876 294652 527882 294704
rect 12434 294584 12440 294636
rect 12492 294624 12498 294636
rect 241882 294624 241888 294636
rect 12492 294596 241888 294624
rect 12492 294584 12498 294596
rect 241882 294584 241888 294596
rect 241940 294584 241946 294636
rect 324958 294584 324964 294636
rect 325016 294624 325022 294636
rect 542354 294624 542360 294636
rect 325016 294596 542360 294624
rect 325016 294584 325022 294596
rect 542354 294584 542360 294596
rect 542412 294584 542418 294636
rect 3326 293904 3332 293956
rect 3384 293944 3390 293956
rect 224218 293944 224224 293956
rect 3384 293916 224224 293944
rect 3384 293904 3390 293916
rect 224218 293904 224224 293916
rect 224276 293904 224282 293956
rect 323394 293292 323400 293344
rect 323452 293332 323458 293344
rect 534718 293332 534724 293344
rect 323452 293304 534724 293332
rect 323452 293292 323458 293304
rect 534718 293292 534724 293304
rect 534776 293292 534782 293344
rect 93854 293224 93860 293276
rect 93912 293264 93918 293276
rect 254210 293264 254216 293276
rect 93912 293236 254216 293264
rect 93912 293224 93918 293236
rect 254210 293224 254216 293236
rect 254268 293224 254274 293276
rect 328914 293224 328920 293276
rect 328972 293264 328978 293276
rect 571334 293264 571340 293276
rect 328972 293236 571340 293264
rect 328972 293224 328978 293236
rect 571334 293224 571340 293236
rect 571392 293224 571398 293276
rect 97994 291864 98000 291916
rect 98052 291904 98058 291916
rect 255866 291904 255872 291916
rect 98052 291876 255872 291904
rect 98052 291864 98058 291876
rect 255866 291864 255872 291876
rect 255924 291864 255930 291916
rect 313918 291864 313924 291916
rect 313976 291904 313982 291916
rect 476758 291904 476764 291916
rect 313976 291876 476764 291904
rect 313976 291864 313982 291876
rect 476758 291864 476764 291876
rect 476816 291864 476822 291916
rect 75914 291796 75920 291848
rect 75972 291836 75978 291848
rect 251174 291836 251180 291848
rect 75972 291808 251180 291836
rect 75972 291796 75978 291808
rect 251174 291796 251180 291808
rect 251232 291796 251238 291848
rect 323302 291796 323308 291848
rect 323360 291836 323366 291848
rect 538858 291836 538864 291848
rect 323360 291808 538864 291836
rect 323360 291796 323366 291808
rect 538858 291796 538864 291808
rect 538916 291796 538922 291848
rect 78674 290504 78680 290556
rect 78732 290544 78738 290556
rect 251542 290544 251548 290556
rect 78732 290516 251548 290544
rect 78732 290504 78738 290516
rect 251542 290504 251548 290516
rect 251600 290504 251606 290556
rect 22094 290436 22100 290488
rect 22152 290476 22158 290488
rect 243078 290476 243084 290488
rect 22152 290448 243084 290476
rect 22152 290436 22158 290448
rect 243078 290436 243084 290448
rect 243136 290436 243142 290488
rect 327534 290436 327540 290488
rect 327592 290476 327598 290488
rect 563698 290476 563704 290488
rect 327592 290448 563704 290476
rect 327592 290436 327598 290448
rect 563698 290436 563704 290448
rect 563756 290436 563762 290488
rect 85574 289144 85580 289196
rect 85632 289184 85638 289196
rect 252830 289184 252836 289196
rect 85632 289156 252836 289184
rect 85632 289144 85638 289156
rect 252830 289144 252836 289156
rect 252888 289144 252894 289196
rect 30374 289076 30380 289128
rect 30432 289116 30438 289128
rect 244826 289116 244832 289128
rect 30432 289088 244832 289116
rect 30432 289076 30438 289088
rect 244826 289076 244832 289088
rect 244884 289076 244890 289128
rect 328822 289076 328828 289128
rect 328880 289116 328886 289128
rect 570598 289116 570604 289128
rect 328880 289088 570604 289116
rect 328880 289076 328886 289088
rect 570598 289076 570604 289088
rect 570656 289076 570662 289128
rect 308214 287716 308220 287768
rect 308272 287756 308278 287768
rect 440326 287756 440332 287768
rect 308272 287728 440332 287756
rect 308272 287716 308278 287728
rect 440326 287716 440332 287728
rect 440384 287716 440390 287768
rect 34514 287648 34520 287700
rect 34572 287688 34578 287700
rect 244550 287688 244556 287700
rect 34572 287660 244556 287688
rect 34572 287648 34578 287660
rect 244550 287648 244556 287660
rect 244608 287648 244614 287700
rect 328730 287648 328736 287700
rect 328788 287688 328794 287700
rect 575474 287688 575480 287700
rect 328788 287660 575480 287688
rect 328788 287648 328794 287660
rect 575474 287648 575480 287660
rect 575532 287648 575538 287700
rect 309502 286424 309508 286476
rect 309560 286464 309566 286476
rect 442350 286464 442356 286476
rect 309560 286436 442356 286464
rect 309560 286424 309566 286436
rect 442350 286424 442356 286436
rect 442408 286424 442414 286476
rect 309594 286356 309600 286408
rect 309652 286396 309658 286408
rect 448514 286396 448520 286408
rect 309652 286368 448520 286396
rect 309652 286356 309658 286368
rect 448514 286356 448520 286368
rect 448572 286356 448578 286408
rect 49694 286288 49700 286340
rect 49752 286328 49758 286340
rect 247402 286328 247408 286340
rect 49752 286300 247408 286328
rect 49752 286288 49758 286300
rect 247402 286288 247408 286300
rect 247460 286288 247466 286340
rect 326246 286288 326252 286340
rect 326304 286328 326310 286340
rect 553394 286328 553400 286340
rect 326304 286300 553400 286328
rect 326304 286288 326310 286300
rect 553394 286288 553400 286300
rect 553452 286288 553458 286340
rect 312538 285064 312544 285116
rect 312596 285104 312602 285116
rect 454034 285104 454040 285116
rect 312596 285076 454040 285104
rect 312596 285064 312602 285076
rect 454034 285064 454040 285076
rect 454092 285064 454098 285116
rect 63494 284996 63500 285048
rect 63552 285036 63558 285048
rect 250070 285036 250076 285048
rect 63552 285008 250076 285036
rect 63552 284996 63558 285008
rect 250070 284996 250076 285008
rect 250128 284996 250134 285048
rect 313826 284996 313832 285048
rect 313884 285036 313890 285048
rect 471238 285036 471244 285048
rect 313884 285008 471244 285036
rect 313884 284996 313890 285008
rect 471238 284996 471244 285008
rect 471296 284996 471302 285048
rect 26234 284928 26240 284980
rect 26292 284968 26298 284980
rect 242986 284968 242992 284980
rect 26292 284940 242992 284968
rect 26292 284928 26298 284940
rect 242986 284928 242992 284940
rect 243044 284928 243050 284980
rect 327442 284928 327448 284980
rect 327500 284968 327506 284980
rect 560938 284968 560944 284980
rect 327500 284940 560944 284968
rect 327500 284928 327506 284940
rect 560938 284928 560944 284940
rect 560996 284928 561002 284980
rect 77294 283636 77300 283688
rect 77352 283676 77358 283688
rect 251450 283676 251456 283688
rect 77352 283648 251456 283676
rect 77352 283636 77358 283648
rect 251450 283636 251456 283648
rect 251508 283636 251514 283688
rect 313642 283636 313648 283688
rect 313700 283676 313706 283688
rect 471974 283676 471980 283688
rect 313700 283648 471980 283676
rect 313700 283636 313706 283648
rect 471974 283636 471980 283648
rect 472032 283636 472038 283688
rect 40034 283568 40040 283620
rect 40092 283608 40098 283620
rect 245930 283608 245936 283620
rect 40092 283580 245936 283608
rect 40092 283568 40098 283580
rect 245930 283568 245936 283580
rect 245988 283568 245994 283620
rect 313734 283568 313740 283620
rect 313792 283608 313798 283620
rect 473446 283608 473452 283620
rect 313792 283580 473452 283608
rect 313792 283568 313798 283580
rect 473446 283568 473452 283580
rect 473504 283568 473510 283620
rect 310882 282276 310888 282328
rect 310940 282316 310946 282328
rect 452654 282316 452660 282328
rect 310940 282288 452660 282316
rect 310940 282276 310946 282288
rect 452654 282276 452660 282288
rect 452712 282276 452718 282328
rect 81434 282208 81440 282260
rect 81492 282248 81498 282260
rect 252738 282248 252744 282260
rect 81492 282220 252744 282248
rect 81492 282208 81498 282220
rect 252738 282208 252744 282220
rect 252796 282208 252802 282260
rect 310790 282208 310796 282260
rect 310848 282248 310854 282260
rect 460934 282248 460940 282260
rect 310848 282220 460940 282248
rect 310848 282208 310854 282220
rect 460934 282208 460940 282220
rect 460992 282208 460998 282260
rect 44174 282140 44180 282192
rect 44232 282180 44238 282192
rect 245838 282180 245844 282192
rect 44232 282152 245844 282180
rect 44232 282140 44238 282152
rect 245838 282140 245844 282152
rect 245896 282140 245902 282192
rect 319162 282140 319168 282192
rect 319220 282180 319226 282192
rect 506566 282180 506572 282192
rect 319220 282152 506572 282180
rect 319220 282140 319226 282152
rect 506566 282140 506572 282152
rect 506624 282140 506630 282192
rect 309410 280848 309416 280900
rect 309468 280888 309474 280900
rect 444374 280888 444380 280900
rect 309468 280860 444380 280888
rect 309468 280848 309474 280860
rect 444374 280848 444380 280860
rect 444432 280848 444438 280900
rect 4890 280780 4896 280832
rect 4948 280820 4954 280832
rect 240318 280820 240324 280832
rect 4948 280792 240324 280820
rect 4948 280780 4954 280792
rect 240318 280780 240324 280792
rect 240376 280780 240382 280832
rect 319070 280780 319076 280832
rect 319128 280820 319134 280832
rect 509234 280820 509240 280832
rect 319128 280792 509240 280820
rect 319128 280780 319134 280792
rect 509234 280780 509240 280792
rect 509292 280780 509298 280832
rect 309318 279488 309324 279540
rect 309376 279528 309382 279540
rect 446398 279528 446404 279540
rect 309376 279500 446404 279528
rect 309376 279488 309382 279500
rect 446398 279488 446404 279500
rect 446456 279488 446462 279540
rect 10410 279420 10416 279472
rect 10468 279460 10474 279472
rect 240502 279460 240508 279472
rect 10468 279432 240508 279460
rect 10468 279420 10474 279432
rect 240502 279420 240508 279432
rect 240560 279420 240566 279472
rect 317690 279420 317696 279472
rect 317748 279460 317754 279472
rect 499574 279460 499580 279472
rect 317748 279432 499580 279460
rect 317748 279420 317754 279432
rect 499574 279420 499580 279432
rect 499632 279420 499638 279472
rect 310698 278060 310704 278112
rect 310756 278100 310762 278112
rect 457438 278100 457444 278112
rect 310756 278072 457444 278100
rect 310756 278060 310762 278072
rect 457438 278060 457444 278072
rect 457496 278060 457502 278112
rect 320450 277992 320456 278044
rect 320508 278032 320514 278044
rect 517514 278032 517520 278044
rect 320508 278004 517520 278032
rect 320508 277992 320514 278004
rect 517514 277992 517520 278004
rect 517572 277992 517578 278044
rect 312262 276700 312268 276752
rect 312320 276740 312326 276752
rect 460198 276740 460204 276752
rect 312320 276712 460204 276740
rect 312320 276700 312326 276712
rect 460198 276700 460204 276712
rect 460256 276700 460262 276752
rect 320358 276632 320364 276684
rect 320416 276672 320422 276684
rect 521654 276672 521660 276684
rect 320416 276644 521660 276672
rect 320416 276632 320422 276644
rect 521654 276632 521660 276644
rect 521712 276632 521718 276684
rect 312170 275340 312176 275392
rect 312228 275380 312234 275392
rect 464338 275380 464344 275392
rect 312228 275352 464344 275380
rect 312228 275340 312234 275352
rect 464338 275340 464344 275352
rect 464396 275340 464402 275392
rect 55214 275272 55220 275324
rect 55272 275312 55278 275324
rect 248690 275312 248696 275324
rect 55272 275284 248696 275312
rect 55272 275272 55278 275284
rect 248690 275272 248696 275284
rect 248748 275272 248754 275324
rect 323210 275272 323216 275324
rect 323268 275312 323274 275324
rect 539686 275312 539692 275324
rect 323268 275284 539692 275312
rect 323268 275272 323274 275284
rect 539686 275272 539692 275284
rect 539744 275272 539750 275324
rect 59354 273912 59360 273964
rect 59412 273952 59418 273964
rect 248598 273952 248604 273964
rect 59412 273924 248604 273952
rect 59412 273912 59418 273924
rect 248598 273912 248604 273924
rect 248656 273912 248662 273964
rect 312078 273912 312084 273964
rect 312136 273952 312142 273964
rect 467098 273952 467104 273964
rect 312136 273924 467104 273952
rect 312136 273912 312142 273924
rect 467098 273912 467104 273924
rect 467156 273912 467162 273964
rect 364978 273164 364984 273216
rect 365036 273204 365042 273216
rect 579890 273204 579896 273216
rect 365036 273176 579896 273204
rect 365036 273164 365042 273176
rect 579890 273164 579896 273176
rect 579948 273164 579954 273216
rect 62114 272484 62120 272536
rect 62172 272524 62178 272536
rect 249978 272524 249984 272536
rect 62172 272496 249984 272524
rect 62172 272484 62178 272496
rect 249978 272484 249984 272496
rect 250036 272484 250042 272536
rect 308122 271328 308128 271380
rect 308180 271368 308186 271380
rect 436738 271368 436744 271380
rect 308180 271340 436744 271368
rect 308180 271328 308186 271340
rect 436738 271328 436744 271340
rect 436796 271328 436802 271380
rect 313550 271260 313556 271312
rect 313608 271300 313614 271312
rect 475378 271300 475384 271312
rect 313608 271272 475384 271300
rect 313608 271260 313614 271272
rect 475378 271260 475384 271272
rect 475436 271260 475442 271312
rect 327350 271192 327356 271244
rect 327408 271232 327414 271244
rect 560294 271232 560300 271244
rect 327408 271204 560300 271232
rect 327408 271192 327414 271204
rect 560294 271192 560300 271204
rect 560352 271192 560358 271244
rect 66254 271124 66260 271176
rect 66312 271164 66318 271176
rect 250346 271164 250352 271176
rect 66312 271136 250352 271164
rect 66312 271124 66318 271136
rect 250346 271124 250352 271136
rect 250404 271124 250410 271176
rect 328638 271124 328644 271176
rect 328696 271164 328702 271176
rect 567838 271164 567844 271176
rect 328696 271136 567844 271164
rect 328696 271124 328702 271136
rect 567838 271124 567844 271136
rect 567896 271124 567902 271176
rect 314930 269968 314936 270020
rect 314988 270008 314994 270020
rect 481634 270008 481640 270020
rect 314988 269980 481640 270008
rect 314988 269968 314994 269980
rect 481634 269968 481640 269980
rect 481692 269968 481698 270020
rect 326154 269900 326160 269952
rect 326212 269940 326218 269952
rect 556154 269940 556160 269952
rect 326212 269912 556160 269940
rect 326212 269900 326218 269912
rect 556154 269900 556160 269912
rect 556212 269900 556218 269952
rect 327258 269832 327264 269884
rect 327316 269872 327322 269884
rect 567194 269872 567200 269884
rect 327316 269844 567200 269872
rect 327316 269832 327322 269844
rect 567194 269832 567200 269844
rect 567252 269832 567258 269884
rect 73154 269764 73160 269816
rect 73212 269804 73218 269816
rect 251358 269804 251364 269816
rect 73212 269776 251364 269804
rect 73212 269764 73218 269776
rect 251358 269764 251364 269776
rect 251416 269764 251422 269816
rect 328546 269764 328552 269816
rect 328604 269804 328610 269816
rect 571978 269804 571984 269816
rect 328604 269776 571984 269804
rect 328604 269764 328610 269776
rect 571978 269764 571984 269776
rect 572036 269764 572042 269816
rect 313366 268676 313372 268728
rect 313424 268716 313430 268728
rect 474734 268716 474740 268728
rect 313424 268688 474740 268716
rect 313424 268676 313430 268688
rect 474734 268676 474740 268688
rect 474792 268676 474798 268728
rect 313458 268608 313464 268660
rect 313516 268648 313522 268660
rect 477494 268648 477500 268660
rect 313516 268620 477500 268648
rect 313516 268608 313522 268620
rect 477494 268608 477500 268620
rect 477552 268608 477558 268660
rect 314838 268540 314844 268592
rect 314896 268580 314902 268592
rect 484394 268580 484400 268592
rect 314896 268552 484400 268580
rect 314896 268540 314902 268552
rect 484394 268540 484400 268552
rect 484452 268540 484458 268592
rect 322198 268472 322204 268524
rect 322256 268512 322262 268524
rect 524414 268512 524420 268524
rect 322256 268484 524420 268512
rect 322256 268472 322262 268484
rect 524414 268472 524420 268484
rect 524472 268472 524478 268524
rect 324774 268404 324780 268456
rect 324832 268444 324838 268456
rect 546494 268444 546500 268456
rect 324832 268416 546500 268444
rect 324832 268404 324838 268416
rect 546494 268404 546500 268416
rect 546552 268404 546558 268456
rect 77386 268336 77392 268388
rect 77444 268376 77450 268388
rect 251726 268376 251732 268388
rect 77444 268348 251732 268376
rect 77444 268336 77450 268348
rect 251726 268336 251732 268348
rect 251784 268336 251790 268388
rect 324866 268336 324872 268388
rect 324924 268376 324930 268388
rect 549254 268376 549260 268388
rect 324924 268348 549260 268376
rect 324924 268336 324930 268348
rect 549254 268336 549260 268348
rect 549312 268336 549318 268388
rect 2958 267656 2964 267708
rect 3016 267696 3022 267708
rect 225598 267696 225604 267708
rect 3016 267668 225604 267696
rect 3016 267656 3022 267668
rect 225598 267656 225604 267668
rect 225656 267656 225662 267708
rect 314746 267112 314752 267164
rect 314804 267152 314810 267164
rect 485774 267152 485780 267164
rect 314804 267124 485780 267152
rect 314804 267112 314810 267124
rect 485774 267112 485780 267124
rect 485832 267112 485838 267164
rect 316494 267044 316500 267096
rect 316552 267084 316558 267096
rect 492674 267084 492680 267096
rect 316552 267056 492680 267084
rect 316552 267044 316558 267056
rect 492674 267044 492680 267056
rect 492732 267044 492738 267096
rect 317598 266976 317604 267028
rect 317656 267016 317662 267028
rect 494790 267016 494796 267028
rect 317656 266988 494796 267016
rect 317656 266976 317662 266988
rect 494790 266976 494796 266988
rect 494848 266976 494854 267028
rect 84194 265684 84200 265736
rect 84252 265724 84258 265736
rect 253014 265724 253020 265736
rect 84252 265696 253020 265724
rect 84252 265684 84258 265696
rect 253014 265684 253020 265696
rect 253072 265684 253078 265736
rect 316402 265684 316408 265736
rect 316460 265724 316466 265736
rect 496814 265724 496820 265736
rect 316460 265696 496820 265724
rect 316460 265684 316466 265696
rect 496814 265684 496820 265696
rect 496872 265684 496878 265736
rect 7650 265616 7656 265668
rect 7708 265656 7714 265668
rect 240410 265656 240416 265668
rect 7708 265628 240416 265656
rect 7708 265616 7714 265628
rect 240410 265616 240416 265628
rect 240468 265616 240474 265668
rect 317506 265616 317512 265668
rect 317564 265656 317570 265668
rect 502334 265656 502340 265668
rect 317564 265628 502340 265656
rect 317564 265616 317570 265628
rect 502334 265616 502340 265628
rect 502392 265616 502398 265668
rect 317414 264324 317420 264376
rect 317472 264364 317478 264376
rect 503714 264364 503720 264376
rect 317472 264336 503720 264364
rect 317472 264324 317478 264336
rect 503714 264324 503720 264336
rect 503772 264324 503778 264376
rect 318978 264256 318984 264308
rect 319036 264296 319042 264308
rect 511258 264296 511264 264308
rect 319036 264268 511264 264296
rect 319036 264256 319042 264268
rect 511258 264256 511264 264268
rect 511316 264256 511322 264308
rect 17954 264188 17960 264240
rect 18012 264228 18018 264240
rect 241790 264228 241796 264240
rect 18012 264200 241796 264228
rect 18012 264188 18018 264200
rect 241790 264188 241796 264200
rect 241848 264188 241854 264240
rect 326062 264188 326068 264240
rect 326120 264228 326126 264240
rect 556246 264228 556252 264240
rect 326120 264200 556252 264228
rect 326120 264188 326126 264200
rect 556246 264188 556252 264200
rect 556304 264188 556310 264240
rect 318886 263100 318892 263152
rect 318944 263140 318950 263152
rect 510614 263140 510620 263152
rect 318944 263112 510620 263140
rect 318944 263100 318950 263112
rect 510614 263100 510620 263112
rect 510672 263100 510678 263152
rect 320266 263032 320272 263084
rect 320324 263072 320330 263084
rect 516134 263072 516140 263084
rect 320324 263044 516140 263072
rect 320324 263032 320330 263044
rect 516134 263032 516140 263044
rect 516192 263032 516198 263084
rect 324682 262964 324688 263016
rect 324740 263004 324746 263016
rect 545114 263004 545120 263016
rect 324740 262976 545120 263004
rect 324740 262964 324746 262976
rect 545114 262964 545120 262976
rect 545172 262964 545178 263016
rect 324590 262896 324596 262948
rect 324648 262936 324654 262948
rect 547874 262936 547880 262948
rect 324648 262908 547880 262936
rect 324648 262896 324654 262908
rect 547874 262896 547880 262908
rect 547932 262896 547938 262948
rect 41414 262828 41420 262880
rect 41472 262868 41478 262880
rect 246114 262868 246120 262880
rect 41472 262840 246120 262868
rect 41472 262828 41478 262840
rect 246114 262828 246120 262840
rect 246172 262828 246178 262880
rect 325970 262828 325976 262880
rect 326028 262868 326034 262880
rect 552014 262868 552020 262880
rect 326028 262840 552020 262868
rect 326028 262828 326034 262840
rect 552014 262828 552020 262840
rect 552072 262828 552078 262880
rect 320174 261672 320180 261724
rect 320232 261712 320238 261724
rect 520274 261712 520280 261724
rect 320232 261684 520280 261712
rect 320232 261672 320238 261684
rect 520274 261672 520280 261684
rect 520332 261672 520338 261724
rect 322106 261604 322112 261656
rect 322164 261644 322170 261656
rect 531314 261644 531320 261656
rect 322164 261616 531320 261644
rect 322164 261604 322170 261616
rect 531314 261604 531320 261616
rect 531372 261604 531378 261656
rect 323118 261536 323124 261588
rect 323176 261576 323182 261588
rect 535454 261576 535460 261588
rect 323176 261548 535460 261576
rect 323176 261536 323182 261548
rect 535454 261536 535460 261548
rect 535512 261536 535518 261588
rect 324498 261468 324504 261520
rect 324556 261508 324562 261520
rect 540974 261508 540980 261520
rect 324556 261480 540980 261508
rect 324556 261468 324562 261480
rect 540974 261468 540980 261480
rect 541032 261468 541038 261520
rect 311986 260312 311992 260364
rect 312044 260352 312050 260364
rect 466454 260352 466460 260364
rect 312044 260324 466460 260352
rect 312044 260312 312050 260324
rect 466454 260312 466460 260324
rect 466512 260312 466518 260364
rect 316310 260244 316316 260296
rect 316368 260284 316374 260296
rect 495434 260284 495440 260296
rect 316368 260256 495440 260284
rect 316368 260244 316374 260256
rect 495434 260244 495440 260256
rect 495492 260244 495498 260296
rect 322014 260176 322020 260228
rect 322072 260216 322078 260228
rect 527174 260216 527180 260228
rect 322072 260188 527180 260216
rect 322072 260176 322078 260188
rect 527174 260176 527180 260188
rect 527232 260176 527238 260228
rect 11698 260108 11704 260160
rect 11756 260148 11762 260160
rect 241698 260148 241704 260160
rect 11756 260120 241704 260148
rect 11756 260108 11762 260120
rect 241698 260108 241704 260120
rect 241756 260108 241762 260160
rect 363598 260108 363604 260160
rect 363656 260148 363662 260160
rect 580442 260148 580448 260160
rect 363656 260120 580448 260148
rect 363656 260108 363662 260120
rect 580442 260108 580448 260120
rect 580500 260108 580506 260160
rect 313274 258884 313280 258936
rect 313332 258924 313338 258936
rect 470594 258924 470600 258936
rect 313332 258896 470600 258924
rect 313332 258884 313338 258896
rect 470594 258884 470600 258896
rect 470652 258884 470658 258936
rect 316126 258816 316132 258868
rect 316184 258856 316190 258868
rect 488534 258856 488540 258868
rect 316184 258828 488540 258856
rect 316184 258816 316190 258828
rect 488534 258816 488540 258828
rect 488592 258816 488598 258868
rect 316218 258748 316224 258800
rect 316276 258788 316282 258800
rect 491294 258788 491300 258800
rect 316276 258760 491300 258788
rect 316276 258748 316282 258760
rect 491294 258748 491300 258760
rect 491352 258748 491358 258800
rect 56594 258680 56600 258732
rect 56652 258720 56658 258732
rect 248966 258720 248972 258732
rect 56652 258692 248972 258720
rect 56652 258680 56658 258692
rect 248966 258680 248972 258692
rect 249024 258680 249030 258732
rect 360838 258680 360844 258732
rect 360896 258720 360902 258732
rect 580350 258720 580356 258732
rect 360896 258692 580356 258720
rect 360896 258680 360902 258692
rect 580350 258680 580356 258692
rect 580408 258680 580414 258732
rect 321922 257320 321928 257372
rect 321980 257360 321986 257372
rect 523126 257360 523132 257372
rect 321980 257332 523132 257360
rect 321980 257320 321986 257332
rect 523126 257320 523132 257332
rect 523184 257320 523190 257372
rect 297910 256096 297916 256148
rect 297968 256136 297974 256148
rect 330110 256136 330116 256148
rect 297968 256108 330116 256136
rect 297968 256096 297974 256108
rect 330110 256096 330116 256108
rect 330168 256096 330174 256148
rect 297634 256028 297640 256080
rect 297692 256068 297698 256080
rect 332686 256068 332692 256080
rect 297692 256040 332692 256068
rect 297692 256028 297698 256040
rect 332686 256028 332692 256040
rect 332744 256028 332750 256080
rect 297266 255960 297272 256012
rect 297324 256000 297330 256012
rect 336918 256000 336924 256012
rect 297324 255972 336924 256000
rect 297324 255960 297330 255972
rect 336918 255960 336924 255972
rect 336976 255960 336982 256012
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 157978 255252 157984 255264
rect 3200 255224 157984 255252
rect 3200 255212 3206 255224
rect 157978 255212 157984 255224
rect 158036 255212 158042 255264
rect 238478 254532 238484 254584
rect 238536 254572 238542 254584
rect 346762 254572 346768 254584
rect 238536 254544 346768 254572
rect 238536 254532 238542 254544
rect 346762 254532 346768 254544
rect 346820 254532 346826 254584
rect 373258 254532 373264 254584
rect 373316 254572 373322 254584
rect 581086 254572 581092 254584
rect 373316 254544 581092 254572
rect 373316 254532 373322 254544
rect 581086 254532 581092 254544
rect 581144 254532 581150 254584
rect 60826 253172 60832 253224
rect 60884 253212 60890 253224
rect 248874 253212 248880 253224
rect 60884 253184 248880 253212
rect 60884 253172 60890 253184
rect 248874 253172 248880 253184
rect 248932 253172 248938 253224
rect 307846 253172 307852 253224
rect 307904 253212 307910 253224
rect 442994 253212 443000 253224
rect 307904 253184 443000 253212
rect 307904 253172 307910 253184
rect 442994 253172 443000 253184
rect 443052 253172 443058 253224
rect 315298 251948 315304 252000
rect 315356 251988 315362 252000
rect 467834 251988 467840 252000
rect 315356 251960 467840 251988
rect 315356 251948 315362 251960
rect 467834 251948 467840 251960
rect 467892 251948 467898 252000
rect 321830 251880 321836 251932
rect 321888 251920 321894 251932
rect 528554 251920 528560 251932
rect 321888 251892 528560 251920
rect 321888 251880 321894 251892
rect 528554 251880 528560 251892
rect 528612 251880 528618 251932
rect 74534 251812 74540 251864
rect 74592 251852 74598 251864
rect 251634 251852 251640 251864
rect 74592 251824 251640 251852
rect 74592 251812 74598 251824
rect 251634 251812 251640 251824
rect 251692 251812 251698 251864
rect 321738 251812 321744 251864
rect 321796 251852 321802 251864
rect 531406 251852 531412 251864
rect 321796 251824 531412 251852
rect 321796 251812 321802 251824
rect 531406 251812 531412 251824
rect 531464 251812 531470 251864
rect 288342 251132 288348 251184
rect 288400 251172 288406 251184
rect 334066 251172 334072 251184
rect 288400 251144 334072 251172
rect 288400 251132 288406 251144
rect 334066 251132 334072 251144
rect 334124 251132 334130 251184
rect 293586 251064 293592 251116
rect 293644 251104 293650 251116
rect 339586 251104 339592 251116
rect 293644 251076 339592 251104
rect 293644 251064 293650 251076
rect 339586 251064 339592 251076
rect 339644 251064 339650 251116
rect 292390 250996 292396 251048
rect 292448 251036 292454 251048
rect 339954 251036 339960 251048
rect 292448 251008 339960 251036
rect 292448 250996 292454 251008
rect 339954 250996 339960 251008
rect 340012 250996 340018 251048
rect 290918 250928 290924 250980
rect 290976 250968 290982 250980
rect 338298 250968 338304 250980
rect 290976 250940 338304 250968
rect 290976 250928 290982 250940
rect 338298 250928 338304 250940
rect 338356 250928 338362 250980
rect 291010 250860 291016 250912
rect 291068 250900 291074 250912
rect 338390 250900 338396 250912
rect 291068 250872 338396 250900
rect 291068 250860 291074 250872
rect 338390 250860 338396 250872
rect 338448 250860 338454 250912
rect 275922 250792 275928 250844
rect 275980 250832 275986 250844
rect 331950 250832 331956 250844
rect 275980 250804 331956 250832
rect 275980 250792 275986 250804
rect 331950 250792 331956 250804
rect 332008 250792 332014 250844
rect 349430 250792 349436 250844
rect 349488 250832 349494 250844
rect 438210 250832 438216 250844
rect 349488 250804 438216 250832
rect 349488 250792 349494 250804
rect 438210 250792 438216 250804
rect 438268 250792 438274 250844
rect 283926 250724 283932 250776
rect 283984 250764 283990 250776
rect 342438 250764 342444 250776
rect 283984 250736 342444 250764
rect 283984 250724 283990 250736
rect 342438 250724 342444 250736
rect 342496 250724 342502 250776
rect 349338 250724 349344 250776
rect 349396 250764 349402 250776
rect 441706 250764 441712 250776
rect 349396 250736 441712 250764
rect 349396 250724 349402 250736
rect 441706 250724 441712 250736
rect 441764 250724 441770 250776
rect 281258 250656 281264 250708
rect 281316 250696 281322 250708
rect 342530 250696 342536 250708
rect 281316 250668 342536 250696
rect 281316 250656 281322 250668
rect 342530 250656 342536 250668
rect 342588 250656 342594 250708
rect 349614 250656 349620 250708
rect 349672 250696 349678 250708
rect 441798 250696 441804 250708
rect 349672 250668 441804 250696
rect 349672 250656 349678 250668
rect 441798 250656 441804 250668
rect 441856 250656 441862 250708
rect 310606 250588 310612 250640
rect 310664 250628 310670 250640
rect 456886 250628 456892 250640
rect 310664 250600 456892 250628
rect 310664 250588 310670 250600
rect 456886 250588 456892 250600
rect 456944 250588 456950 250640
rect 310514 250520 310520 250572
rect 310572 250560 310578 250572
rect 459554 250560 459560 250572
rect 310572 250532 459560 250560
rect 310572 250520 310578 250532
rect 459554 250520 459560 250532
rect 459612 250520 459618 250572
rect 13814 250452 13820 250504
rect 13872 250492 13878 250504
rect 242066 250492 242072 250504
rect 13872 250464 242072 250492
rect 13872 250452 13878 250464
rect 242066 250452 242072 250464
rect 242124 250452 242130 250504
rect 318794 250452 318800 250504
rect 318852 250492 318858 250504
rect 514110 250492 514116 250504
rect 318852 250464 514116 250492
rect 318852 250452 318858 250464
rect 514110 250452 514116 250464
rect 514168 250452 514174 250504
rect 296438 250384 296444 250436
rect 296496 250424 296502 250436
rect 341150 250424 341156 250436
rect 296496 250396 341156 250424
rect 296496 250384 296502 250396
rect 341150 250384 341156 250396
rect 341208 250384 341214 250436
rect 289630 250316 289636 250368
rect 289688 250356 289694 250368
rect 334158 250356 334164 250368
rect 289688 250328 334164 250356
rect 289688 250316 289694 250328
rect 334158 250316 334164 250328
rect 334216 250316 334222 250368
rect 299290 250248 299296 250300
rect 299348 250288 299354 250300
rect 341058 250288 341064 250300
rect 299348 250260 341064 250288
rect 299348 250248 299354 250260
rect 341058 250248 341064 250260
rect 341116 250248 341122 250300
rect 296898 249432 296904 249484
rect 296956 249472 296962 249484
rect 297358 249472 297364 249484
rect 296956 249444 297364 249472
rect 296956 249432 296962 249444
rect 297358 249432 297364 249444
rect 297416 249432 297422 249484
rect 309226 249228 309232 249280
rect 309284 249268 309290 249280
rect 445754 249268 445760 249280
rect 309284 249240 445760 249268
rect 309284 249228 309290 249240
rect 445754 249228 445760 249240
rect 445812 249228 445818 249280
rect 314654 249160 314660 249212
rect 314712 249200 314718 249212
rect 481726 249200 481732 249212
rect 314712 249172 481732 249200
rect 314712 249160 314718 249172
rect 481726 249160 481732 249172
rect 481784 249160 481790 249212
rect 297174 249092 297180 249144
rect 297232 249092 297238 249144
rect 325878 249092 325884 249144
rect 325936 249132 325942 249144
rect 554774 249132 554780 249144
rect 325936 249104 554780 249132
rect 325936 249092 325942 249104
rect 554774 249092 554780 249104
rect 554832 249092 554838 249144
rect 297192 248872 297220 249092
rect 325786 249024 325792 249076
rect 325844 249064 325850 249076
rect 557534 249064 557540 249076
rect 325844 249036 557540 249064
rect 325844 249024 325850 249036
rect 557534 249024 557540 249036
rect 557592 249024 557598 249076
rect 297174 248820 297180 248872
rect 297232 248820 297238 248872
rect 293402 248344 293408 248396
rect 293460 248384 293466 248396
rect 303982 248384 303988 248396
rect 293460 248356 303988 248384
rect 293460 248344 293466 248356
rect 303982 248344 303988 248356
rect 304040 248344 304046 248396
rect 298830 248276 298836 248328
rect 298888 248316 298894 248328
rect 348234 248316 348240 248328
rect 298888 248288 348240 248316
rect 298888 248276 298894 248288
rect 348234 248276 348240 248288
rect 348292 248276 348298 248328
rect 282546 248208 282552 248260
rect 282604 248248 282610 248260
rect 337194 248248 337200 248260
rect 282604 248220 337200 248248
rect 282604 248208 282610 248220
rect 337194 248208 337200 248220
rect 337252 248208 337258 248260
rect 346486 248208 346492 248260
rect 346544 248248 346550 248260
rect 436922 248248 436928 248260
rect 346544 248220 436928 248248
rect 346544 248208 346550 248220
rect 436922 248208 436928 248220
rect 436980 248208 436986 248260
rect 278590 248140 278596 248192
rect 278648 248180 278654 248192
rect 341426 248180 341432 248192
rect 278648 248152 341432 248180
rect 278648 248140 278654 248152
rect 341426 248140 341432 248152
rect 341484 248140 341490 248192
rect 346670 248140 346676 248192
rect 346728 248180 346734 248192
rect 438302 248180 438308 248192
rect 346728 248152 438308 248180
rect 346728 248140 346734 248152
rect 438302 248140 438308 248152
rect 438360 248140 438366 248192
rect 278682 248072 278688 248124
rect 278740 248112 278746 248124
rect 346578 248112 346584 248124
rect 278740 248084 346584 248112
rect 278740 248072 278746 248084
rect 346578 248072 346584 248084
rect 346636 248072 346642 248124
rect 347958 248072 347964 248124
rect 348016 248112 348022 248124
rect 441890 248112 441896 248124
rect 348016 248084 441896 248112
rect 348016 248072 348022 248084
rect 441890 248072 441896 248084
rect 441948 248072 441954 248124
rect 283926 248004 283932 248056
rect 283984 248044 283990 248056
rect 304166 248044 304172 248056
rect 283984 248016 304172 248044
rect 283984 248004 283990 248016
rect 304166 248004 304172 248016
rect 304224 248004 304230 248056
rect 305546 248004 305552 248056
rect 305604 248044 305610 248056
rect 437474 248044 437480 248056
rect 305604 248016 437480 248044
rect 305604 248004 305610 248016
rect 437474 248004 437480 248016
rect 437532 248004 437538 248056
rect 286594 247936 286600 247988
rect 286652 247976 286658 247988
rect 302878 247976 302884 247988
rect 286652 247948 302884 247976
rect 286652 247936 286658 247948
rect 302878 247936 302884 247948
rect 302936 247936 302942 247988
rect 305362 247936 305368 247988
rect 305420 247976 305426 247988
rect 437566 247976 437572 247988
rect 305420 247948 437572 247976
rect 305420 247936 305426 247948
rect 437566 247936 437572 247948
rect 437624 247936 437630 247988
rect 287790 247868 287796 247920
rect 287848 247908 287854 247920
rect 302602 247908 302608 247920
rect 287848 247880 302608 247908
rect 287848 247868 287854 247880
rect 302602 247868 302608 247880
rect 302660 247868 302666 247920
rect 306926 247868 306932 247920
rect 306984 247908 306990 247920
rect 440418 247908 440424 247920
rect 306984 247880 440424 247908
rect 306984 247868 306990 247880
rect 440418 247868 440424 247880
rect 440476 247868 440482 247920
rect 289170 247800 289176 247852
rect 289228 247840 289234 247852
rect 302786 247840 302792 247852
rect 289228 247812 302792 247840
rect 289228 247800 289234 247812
rect 302786 247800 302792 247812
rect 302844 247800 302850 247852
rect 305454 247800 305460 247852
rect 305512 247840 305518 247852
rect 438946 247840 438952 247852
rect 305512 247812 438952 247840
rect 305512 247800 305518 247812
rect 438946 247800 438952 247812
rect 439004 247800 439010 247852
rect 285030 247732 285036 247784
rect 285088 247772 285094 247784
rect 302694 247772 302700 247784
rect 285088 247744 302700 247772
rect 285088 247732 285094 247744
rect 302694 247732 302700 247744
rect 302752 247732 302758 247784
rect 306834 247732 306840 247784
rect 306892 247772 306898 247784
rect 440510 247772 440516 247784
rect 306892 247744 440516 247772
rect 306892 247732 306898 247744
rect 440510 247732 440516 247744
rect 440568 247732 440574 247784
rect 31754 247664 31760 247716
rect 31812 247704 31818 247716
rect 243722 247704 243728 247716
rect 31812 247676 243728 247704
rect 31812 247664 31818 247676
rect 243722 247664 243728 247676
rect 243780 247664 243786 247716
rect 304074 247664 304080 247716
rect 304132 247704 304138 247716
rect 439038 247704 439044 247716
rect 304132 247676 439044 247704
rect 304132 247664 304138 247676
rect 439038 247664 439044 247676
rect 439096 247664 439102 247716
rect 296346 247596 296352 247648
rect 296404 247636 296410 247648
rect 342346 247636 342352 247648
rect 296404 247608 342352 247636
rect 296404 247596 296410 247608
rect 342346 247596 342352 247608
rect 342404 247596 342410 247648
rect 293494 247528 293500 247580
rect 293552 247568 293558 247580
rect 338574 247568 338580 247580
rect 293552 247540 338580 247568
rect 293552 247528 293558 247540
rect 338574 247528 338580 247540
rect 338632 247528 338638 247580
rect 297266 247460 297272 247512
rect 297324 247500 297330 247512
rect 334342 247500 334348 247512
rect 297324 247472 334348 247500
rect 297324 247460 297330 247472
rect 334342 247460 334348 247472
rect 334400 247460 334406 247512
rect 288250 247392 288256 247444
rect 288308 247432 288314 247444
rect 335630 247432 335636 247444
rect 288308 247404 335636 247432
rect 288308 247392 288314 247404
rect 335630 247392 335636 247404
rect 335688 247392 335694 247444
rect 295058 247052 295064 247104
rect 295116 247092 295122 247104
rect 298554 247092 298560 247104
rect 295116 247064 298560 247092
rect 295116 247052 295122 247064
rect 298554 247052 298560 247064
rect 298612 247052 298618 247104
rect 295150 246984 295156 247036
rect 295208 247024 295214 247036
rect 349522 247024 349528 247036
rect 295208 246996 349528 247024
rect 295208 246984 295214 246996
rect 349522 246984 349528 246996
rect 349580 246984 349586 247036
rect 277026 246916 277032 246968
rect 277084 246956 277090 246968
rect 331858 246956 331864 246968
rect 277084 246928 331864 246956
rect 277084 246916 277090 246928
rect 331858 246916 331864 246928
rect 331916 246916 331922 246968
rect 281350 246848 281356 246900
rect 281408 246888 281414 246900
rect 343726 246888 343732 246900
rect 281408 246860 343732 246888
rect 281408 246848 281414 246860
rect 343726 246848 343732 246860
rect 343784 246848 343790 246900
rect 275830 246780 275836 246832
rect 275888 246820 275894 246832
rect 344094 246820 344100 246832
rect 275888 246792 344100 246820
rect 275888 246780 275894 246792
rect 344094 246780 344100 246792
rect 344152 246780 344158 246832
rect 274266 246712 274272 246764
rect 274324 246752 274330 246764
rect 345474 246752 345480 246764
rect 274324 246724 345480 246752
rect 274324 246712 274330 246724
rect 345474 246712 345480 246724
rect 345532 246712 345538 246764
rect 273162 246644 273168 246696
rect 273220 246684 273226 246696
rect 348142 246684 348148 246696
rect 273220 246656 348148 246684
rect 273220 246644 273226 246656
rect 348142 246644 348148 246656
rect 348200 246644 348206 246696
rect 350626 246644 350632 246696
rect 350684 246684 350690 246696
rect 439682 246684 439688 246696
rect 350684 246656 439688 246684
rect 350684 246644 350690 246656
rect 439682 246644 439688 246656
rect 439740 246644 439746 246696
rect 309134 246576 309140 246628
rect 309192 246616 309198 246628
rect 448606 246616 448612 246628
rect 309192 246588 448612 246616
rect 309192 246576 309198 246588
rect 448606 246576 448612 246588
rect 448664 246576 448670 246628
rect 316034 246508 316040 246560
rect 316092 246548 316098 246560
rect 490006 246548 490012 246560
rect 316092 246520 490012 246548
rect 316092 246508 316098 246520
rect 490006 246508 490012 246520
rect 490064 246508 490070 246560
rect 322934 246440 322940 246492
rect 322992 246480 322998 246492
rect 538214 246480 538220 246492
rect 322992 246452 538220 246480
rect 322992 246440 322998 246452
rect 538214 246440 538220 246452
rect 538272 246440 538278 246492
rect 324314 246372 324320 246424
rect 324372 246412 324378 246424
rect 543734 246412 543740 246424
rect 324372 246384 543740 246412
rect 324372 246372 324378 246384
rect 543734 246372 543740 246384
rect 543792 246372 543798 246424
rect 95234 246304 95240 246356
rect 95292 246344 95298 246356
rect 243630 246344 243636 246356
rect 95292 246316 243636 246344
rect 95292 246304 95298 246316
rect 243630 246304 243636 246316
rect 243688 246304 243694 246356
rect 285582 246304 285588 246356
rect 285640 246344 285646 246356
rect 292942 246344 292948 246356
rect 285640 246316 292948 246344
rect 285640 246304 285646 246316
rect 292942 246304 292948 246316
rect 293000 246304 293006 246356
rect 327166 246304 327172 246356
rect 327224 246344 327230 246356
rect 564526 246344 564532 246356
rect 327224 246316 564532 246344
rect 327224 246304 327230 246316
rect 564526 246304 564532 246316
rect 564584 246304 564590 246356
rect 298002 246236 298008 246288
rect 298060 246276 298066 246288
rect 346946 246276 346952 246288
rect 298060 246248 346952 246276
rect 298060 246236 298066 246248
rect 346946 246236 346952 246248
rect 347004 246236 347010 246288
rect 297450 246168 297456 246220
rect 297508 246208 297514 246220
rect 335998 246208 336004 246220
rect 297508 246180 336004 246208
rect 297508 246168 297514 246180
rect 335998 246168 336004 246180
rect 336056 246168 336062 246220
rect 299014 246100 299020 246152
rect 299072 246140 299078 246152
rect 335814 246140 335820 246152
rect 299072 246112 335820 246140
rect 299072 246100 299078 246112
rect 335814 246100 335820 246112
rect 335872 246100 335878 246152
rect 296806 245556 296812 245608
rect 296864 245596 296870 245608
rect 298738 245596 298744 245608
rect 296864 245568 298744 245596
rect 296864 245556 296870 245568
rect 298738 245556 298744 245568
rect 298796 245556 298802 245608
rect 306742 245556 306748 245608
rect 306800 245596 306806 245608
rect 437750 245596 437756 245608
rect 306800 245568 437756 245596
rect 306800 245556 306806 245568
rect 437750 245556 437756 245568
rect 437808 245556 437814 245608
rect 295242 245488 295248 245540
rect 295300 245528 295306 245540
rect 302326 245528 302332 245540
rect 295300 245500 302332 245528
rect 295300 245488 295306 245500
rect 302326 245488 302332 245500
rect 302384 245488 302390 245540
rect 306466 245488 306472 245540
rect 306524 245528 306530 245540
rect 437842 245528 437848 245540
rect 306524 245500 437848 245528
rect 306524 245488 306530 245500
rect 437842 245488 437848 245500
rect 437900 245488 437906 245540
rect 290826 245420 290832 245472
rect 290884 245460 290890 245472
rect 303706 245460 303712 245472
rect 290884 245432 303712 245460
rect 290884 245420 290890 245432
rect 303706 245420 303712 245432
rect 303764 245420 303770 245472
rect 305086 245420 305092 245472
rect 305144 245460 305150 245472
rect 437658 245460 437664 245472
rect 305144 245432 437664 245460
rect 305144 245420 305150 245432
rect 437658 245420 437664 245432
rect 437716 245420 437722 245472
rect 292114 245352 292120 245404
rect 292172 245392 292178 245404
rect 302418 245392 302424 245404
rect 292172 245364 302424 245392
rect 292172 245352 292178 245364
rect 302418 245352 302424 245364
rect 302476 245352 302482 245404
rect 306650 245352 306656 245404
rect 306708 245392 306714 245404
rect 439314 245392 439320 245404
rect 306708 245364 439320 245392
rect 306708 245352 306714 245364
rect 439314 245352 439320 245364
rect 439372 245352 439378 245404
rect 293770 245284 293776 245336
rect 293828 245324 293834 245336
rect 301038 245324 301044 245336
rect 293828 245296 301044 245324
rect 293828 245284 293834 245296
rect 301038 245284 301044 245296
rect 301096 245284 301102 245336
rect 306558 245284 306564 245336
rect 306616 245324 306622 245336
rect 439406 245324 439412 245336
rect 306616 245296 439412 245324
rect 306616 245284 306622 245296
rect 439406 245284 439412 245296
rect 439464 245284 439470 245336
rect 304994 245216 305000 245268
rect 305052 245256 305058 245268
rect 437934 245256 437940 245268
rect 305052 245228 437940 245256
rect 305052 245216 305058 245228
rect 437934 245216 437940 245228
rect 437992 245216 437998 245268
rect 296622 245148 296628 245200
rect 296680 245188 296686 245200
rect 303614 245188 303620 245200
rect 296680 245160 303620 245188
rect 296680 245148 296686 245160
rect 303614 245148 303620 245160
rect 303672 245148 303678 245200
rect 305270 245148 305276 245200
rect 305328 245188 305334 245200
rect 439130 245188 439136 245200
rect 305328 245160 439136 245188
rect 305328 245148 305334 245160
rect 439130 245148 439136 245160
rect 439188 245148 439194 245200
rect 305178 245080 305184 245132
rect 305236 245120 305242 245132
rect 439222 245120 439228 245132
rect 305236 245092 439228 245120
rect 305236 245080 305242 245092
rect 439222 245080 439228 245092
rect 439280 245080 439286 245132
rect 291102 245012 291108 245064
rect 291160 245052 291166 245064
rect 302234 245052 302240 245064
rect 291160 245024 302240 245052
rect 291160 245012 291166 245024
rect 302234 245012 302240 245024
rect 302292 245012 302298 245064
rect 311894 245012 311900 245064
rect 311952 245052 311958 245064
rect 463694 245052 463700 245064
rect 311952 245024 463700 245052
rect 311952 245012 311958 245024
rect 463694 245012 463700 245024
rect 463752 245012 463758 245064
rect 321554 244944 321560 244996
rect 321612 244984 321618 244996
rect 525794 244984 525800 244996
rect 321612 244956 525800 244984
rect 321612 244944 321618 244956
rect 525794 244944 525800 244956
rect 525852 244944 525858 244996
rect 3602 244876 3608 244928
rect 3660 244916 3666 244928
rect 229738 244916 229744 244928
rect 3660 244888 229744 244916
rect 3660 244876 3666 244888
rect 229738 244876 229744 244888
rect 229796 244876 229802 244928
rect 293402 244876 293408 244928
rect 293460 244916 293466 244928
rect 300854 244916 300860 244928
rect 293460 244888 300860 244916
rect 293460 244876 293466 244888
rect 300854 244876 300860 244888
rect 300912 244876 300918 244928
rect 329926 244876 329932 244928
rect 329984 244916 329990 244928
rect 576854 244916 576860 244928
rect 329984 244888 576860 244916
rect 329984 244876 329990 244888
rect 576854 244876 576860 244888
rect 576912 244876 576918 244928
rect 279878 244808 279884 244860
rect 279936 244848 279942 244860
rect 345566 244848 345572 244860
rect 279936 244820 345572 244848
rect 279936 244808 279942 244820
rect 345566 244808 345572 244820
rect 345624 244808 345630 244860
rect 297542 244740 297548 244792
rect 297600 244780 297606 244792
rect 337102 244780 337108 244792
rect 297600 244752 337108 244780
rect 297600 244740 297606 244752
rect 337102 244740 337108 244752
rect 337160 244740 337166 244792
rect 299106 244672 299112 244724
rect 299164 244712 299170 244724
rect 332962 244712 332968 244724
rect 299164 244684 332968 244712
rect 299164 244672 299170 244684
rect 332962 244672 332968 244684
rect 333020 244672 333026 244724
rect 288158 244604 288164 244656
rect 288216 244644 288222 244656
rect 288216 244616 292574 244644
rect 288216 244604 288222 244616
rect 292546 244440 292574 244616
rect 295242 244604 295248 244656
rect 295300 244644 295306 244656
rect 299842 244644 299848 244656
rect 295300 244616 299848 244644
rect 295300 244604 295306 244616
rect 299842 244604 299848 244616
rect 299900 244604 299906 244656
rect 297726 244536 297732 244588
rect 297784 244576 297790 244588
rect 330202 244576 330208 244588
rect 297784 244548 330208 244576
rect 297784 244536 297790 244548
rect 330202 244536 330208 244548
rect 330260 244536 330266 244588
rect 293862 244468 293868 244520
rect 293920 244508 293926 244520
rect 300946 244508 300952 244520
rect 293920 244480 300952 244508
rect 293920 244468 293926 244480
rect 300946 244468 300952 244480
rect 301004 244468 301010 244520
rect 301130 244440 301136 244452
rect 292546 244412 301136 244440
rect 301130 244400 301136 244412
rect 301188 244400 301194 244452
rect 291746 244332 291752 244384
rect 291804 244372 291810 244384
rect 297358 244372 297364 244384
rect 291804 244344 297364 244372
rect 291804 244332 291810 244344
rect 297358 244332 297364 244344
rect 297416 244332 297422 244384
rect 297818 243788 297824 243840
rect 297876 243828 297882 243840
rect 316770 243828 316776 243840
rect 297876 243800 316776 243828
rect 297876 243788 297882 243800
rect 316770 243788 316776 243800
rect 316828 243788 316834 243840
rect 299198 243720 299204 243772
rect 299256 243760 299262 243772
rect 338482 243760 338488 243772
rect 299256 243732 338488 243760
rect 299256 243720 299262 243732
rect 338482 243720 338488 243732
rect 338540 243720 338546 243772
rect 290826 243652 290832 243704
rect 290884 243692 290890 243704
rect 335722 243692 335728 243704
rect 290884 243664 335728 243692
rect 290884 243652 290890 243664
rect 335722 243652 335728 243664
rect 335780 243652 335786 243704
rect 294966 243584 294972 243636
rect 295024 243624 295030 243636
rect 342622 243624 342628 243636
rect 295024 243596 342628 243624
rect 295024 243584 295030 243596
rect 342622 243584 342628 243596
rect 342680 243584 342686 243636
rect 286778 243516 286784 243568
rect 286836 243556 286842 243568
rect 341242 243556 341248 243568
rect 286836 243528 341248 243556
rect 286836 243516 286842 243528
rect 341242 243516 341248 243528
rect 341300 243516 341306 243568
rect 97718 243448 97724 243500
rect 97776 243488 97782 243500
rect 297082 243488 297088 243500
rect 97776 243460 297088 243488
rect 97776 243448 97782 243460
rect 297082 243448 297088 243460
rect 297140 243448 297146 243500
rect 97810 243380 97816 243432
rect 97868 243420 97874 243432
rect 297358 243420 297364 243432
rect 97868 243392 297364 243420
rect 97868 243380 97874 243392
rect 297358 243380 297364 243392
rect 297416 243420 297422 243432
rect 297542 243420 297548 243432
rect 297416 243392 297548 243420
rect 297416 243380 297422 243392
rect 297542 243380 297548 243392
rect 297600 243380 297606 243432
rect 3234 241408 3240 241460
rect 3292 241448 3298 241460
rect 97258 241448 97264 241460
rect 3292 241420 97264 241448
rect 3292 241408 3298 241420
rect 97258 241408 97264 241420
rect 97316 241408 97322 241460
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 95970 215268 95976 215280
rect 3384 215240 95976 215268
rect 3384 215228 3390 215240
rect 95970 215228 95976 215240
rect 96028 215228 96034 215280
rect 3142 188980 3148 189032
rect 3200 189020 3206 189032
rect 94498 189020 94504 189032
rect 3200 188992 94504 189020
rect 3200 188980 3206 188992
rect 94498 188980 94504 188992
rect 94556 188980 94562 189032
rect 3510 164160 3516 164212
rect 3568 164200 3574 164212
rect 93118 164200 93124 164212
rect 3568 164172 93124 164200
rect 3568 164160 3574 164172
rect 93118 164160 93124 164172
rect 93176 164160 93182 164212
rect 297266 243108 297272 243160
rect 297324 243148 297330 243160
rect 297542 243148 297548 243160
rect 297324 243120 297548 243148
rect 297324 243108 297330 243120
rect 297542 243108 297548 243120
rect 297600 243108 297606 243160
rect 293494 239776 293500 239828
rect 293552 239816 293558 239828
rect 293770 239816 293776 239828
rect 293552 239788 293776 239816
rect 293552 239776 293558 239788
rect 293770 239776 293776 239788
rect 293828 239776 293834 239828
rect 297174 195984 297180 196036
rect 297232 196024 297238 196036
rect 298830 196024 298836 196036
rect 297232 195996 298836 196024
rect 297232 195984 297238 195996
rect 298830 195984 298836 195996
rect 298888 195984 298894 196036
rect 295150 195916 295156 195968
rect 295208 195956 295214 195968
rect 297266 195956 297272 195968
rect 295208 195928 297272 195956
rect 295208 195916 295214 195928
rect 297266 195916 297272 195928
rect 297324 195916 297330 195968
rect 280982 193808 280988 193860
rect 281040 193848 281046 193860
rect 297450 193848 297456 193860
rect 281040 193820 297456 193848
rect 281040 193808 281046 193820
rect 297450 193808 297456 193820
rect 297508 193808 297514 193860
rect 283558 191836 283564 191888
rect 283616 191876 283622 191888
rect 299014 191876 299020 191888
rect 283616 191848 299020 191876
rect 283616 191836 283622 191848
rect 299014 191836 299020 191848
rect 299072 191836 299078 191888
rect 297266 189864 297272 189916
rect 297324 189904 297330 189916
rect 298370 189904 298376 189916
rect 297324 189876 298376 189904
rect 297324 189864 297330 189876
rect 298370 189864 298376 189876
rect 298428 189864 298434 189916
rect 238110 174632 238116 174684
rect 238168 174672 238174 174684
rect 260006 174672 260012 174684
rect 238168 174644 260012 174672
rect 238168 174632 238174 174644
rect 260006 174632 260012 174644
rect 260064 174632 260070 174684
rect 245746 174564 245752 174616
rect 245804 174604 245810 174616
rect 277946 174604 277952 174616
rect 245804 174576 277952 174604
rect 245804 174564 245810 174576
rect 277946 174564 277952 174576
rect 278004 174564 278010 174616
rect 237374 174496 237380 174548
rect 237432 174536 237438 174548
rect 276474 174536 276480 174548
rect 237432 174508 276480 174536
rect 237432 174496 237438 174508
rect 276474 174496 276480 174508
rect 276532 174496 276538 174548
rect 239398 173136 239404 173188
rect 239456 173176 239462 173188
rect 266814 173176 266820 173188
rect 239456 173148 266820 173176
rect 239456 173136 239462 173148
rect 266814 173136 266820 173148
rect 266872 173136 266878 173188
rect 282638 171028 282644 171080
rect 282696 171068 282702 171080
rect 297634 171068 297640 171080
rect 282696 171040 297640 171068
rect 282696 171028 282702 171040
rect 297634 171028 297640 171040
rect 297692 171028 297698 171080
rect 297174 170552 297180 170604
rect 297232 170592 297238 170604
rect 298554 170592 298560 170604
rect 297232 170564 298560 170592
rect 297232 170552 297238 170564
rect 298554 170552 298560 170564
rect 298612 170552 298618 170604
rect 238386 170348 238392 170400
rect 238444 170388 238450 170400
rect 282638 170388 282644 170400
rect 238444 170360 282644 170388
rect 238444 170348 238450 170360
rect 282638 170348 282644 170360
rect 282696 170348 282702 170400
rect 293770 168308 293776 168360
rect 293828 168348 293834 168360
rect 297634 168348 297640 168360
rect 293828 168320 297640 168348
rect 293828 168308 293834 168320
rect 297634 168308 297640 168320
rect 297692 168308 297698 168360
rect 238570 167628 238576 167680
rect 238628 167668 238634 167680
rect 297910 167668 297916 167680
rect 238628 167640 297916 167668
rect 238628 167628 238634 167640
rect 297910 167628 297916 167640
rect 297968 167628 297974 167680
rect 97442 159876 97448 159928
rect 97500 159916 97506 159928
rect 297542 159916 297548 159928
rect 97500 159888 297548 159916
rect 97500 159876 97506 159888
rect 297542 159876 297548 159888
rect 297600 159876 297606 159928
rect 97534 159808 97540 159860
rect 97592 159848 97598 159860
rect 297450 159848 297456 159860
rect 97592 159820 297456 159848
rect 97592 159808 97598 159820
rect 297450 159808 297456 159820
rect 297508 159808 297514 159860
rect 97718 159740 97724 159792
rect 97776 159780 97782 159792
rect 283558 159780 283564 159792
rect 97776 159752 283564 159780
rect 97776 159740 97782 159752
rect 283558 159740 283564 159752
rect 283616 159740 283622 159792
rect 97810 159672 97816 159724
rect 97868 159712 97874 159724
rect 280982 159712 280988 159724
rect 97868 159684 280988 159712
rect 97868 159672 97874 159684
rect 280982 159672 280988 159684
rect 281040 159672 281046 159724
rect 97902 159604 97908 159656
rect 97960 159644 97966 159656
rect 238570 159644 238576 159656
rect 97960 159616 238576 159644
rect 97960 159604 97966 159616
rect 238570 159604 238576 159616
rect 238628 159604 238634 159656
rect 286134 159604 286140 159656
rect 286192 159644 286198 159656
rect 299474 159644 299480 159656
rect 286192 159616 299480 159644
rect 286192 159604 286198 159616
rect 299474 159604 299480 159616
rect 299532 159604 299538 159656
rect 97350 159536 97356 159588
rect 97408 159576 97414 159588
rect 238386 159576 238392 159588
rect 97408 159548 238392 159576
rect 97408 159536 97414 159548
rect 238386 159536 238392 159548
rect 238444 159536 238450 159588
rect 287514 159536 287520 159588
rect 287572 159576 287578 159588
rect 302234 159576 302240 159588
rect 287572 159548 302240 159576
rect 287572 159536 287578 159548
rect 302234 159536 302240 159548
rect 302292 159536 302298 159588
rect 288250 159468 288256 159520
rect 288308 159508 288314 159520
rect 335998 159508 336004 159520
rect 288308 159480 336004 159508
rect 288308 159468 288314 159480
rect 335998 159468 336004 159480
rect 336056 159468 336062 159520
rect 289630 159400 289636 159452
rect 289688 159440 289694 159452
rect 338482 159440 338488 159452
rect 289688 159412 338488 159440
rect 289688 159400 289694 159412
rect 338482 159400 338488 159412
rect 338540 159400 338546 159452
rect 173434 159332 173440 159384
rect 173492 159372 173498 159384
rect 294690 159372 294696 159384
rect 173492 159344 294696 159372
rect 173492 159332 173498 159344
rect 294690 159332 294696 159344
rect 294748 159332 294754 159384
rect 297634 159332 297640 159384
rect 297692 159372 297698 159384
rect 348234 159372 348240 159384
rect 297692 159344 348240 159372
rect 297692 159332 297698 159344
rect 348234 159332 348240 159344
rect 348292 159332 348298 159384
rect 291010 159264 291016 159316
rect 291068 159304 291074 159316
rect 350994 159304 351000 159316
rect 291068 159276 351000 159304
rect 291068 159264 291074 159276
rect 350994 159264 351000 159276
rect 351052 159264 351058 159316
rect 290918 159196 290924 159248
rect 290976 159236 290982 159248
rect 353570 159236 353576 159248
rect 290976 159208 353576 159236
rect 290976 159196 290982 159208
rect 353570 159196 353576 159208
rect 353628 159196 353634 159248
rect 206002 159128 206008 159180
rect 206060 159168 206066 159180
rect 267090 159168 267096 159180
rect 206060 159140 267096 159168
rect 206060 159128 206066 159140
rect 267090 159128 267096 159140
rect 267148 159128 267154 159180
rect 293586 159128 293592 159180
rect 293644 159168 293650 159180
rect 356054 159168 356060 159180
rect 293644 159140 356060 159168
rect 293644 159128 293650 159140
rect 356054 159128 356060 159140
rect 356112 159128 356118 159180
rect 165982 159060 165988 159112
rect 166040 159100 166046 159112
rect 238202 159100 238208 159112
rect 166040 159072 238208 159100
rect 166040 159060 166046 159072
rect 238202 159060 238208 159072
rect 238260 159060 238266 159112
rect 299290 159060 299296 159112
rect 299348 159100 299354 159112
rect 363506 159100 363512 159112
rect 299348 159072 363512 159100
rect 299348 159060 299354 159072
rect 363506 159060 363512 159072
rect 363564 159060 363570 159112
rect 156046 158992 156052 159044
rect 156104 159032 156110 159044
rect 243538 159032 243544 159044
rect 156104 159004 243544 159032
rect 156104 158992 156110 159004
rect 243538 158992 243544 159004
rect 243596 158992 243602 159044
rect 296438 158992 296444 159044
rect 296496 159032 296502 159044
rect 360930 159032 360936 159044
rect 296496 159004 360936 159032
rect 296496 158992 296502 159004
rect 360930 158992 360936 159004
rect 360988 158992 360994 159044
rect 158530 158924 158536 158976
rect 158588 158964 158594 158976
rect 257522 158964 257528 158976
rect 158588 158936 257528 158964
rect 158588 158924 158594 158936
rect 257522 158924 257528 158936
rect 257580 158924 257586 158976
rect 281258 158924 281264 158976
rect 281316 158964 281322 158976
rect 370958 158964 370964 158976
rect 281316 158936 370964 158964
rect 281316 158924 281322 158936
rect 370958 158924 370964 158936
rect 371016 158924 371022 158976
rect 284018 158856 284024 158908
rect 284076 158896 284082 158908
rect 368198 158896 368204 158908
rect 284076 158868 368204 158896
rect 284076 158856 284082 158868
rect 368198 158856 368204 158868
rect 368256 158856 368262 158908
rect 168282 158788 168288 158840
rect 168340 158828 168346 158840
rect 284938 158828 284944 158840
rect 168340 158800 284944 158828
rect 168340 158788 168346 158800
rect 284938 158788 284944 158800
rect 284996 158788 285002 158840
rect 292390 158788 292396 158840
rect 292448 158828 292454 158840
rect 358446 158828 358452 158840
rect 292448 158800 358452 158828
rect 292448 158788 292454 158800
rect 358446 158788 358452 158800
rect 358504 158788 358510 158840
rect 160922 158720 160928 158772
rect 160980 158760 160986 158772
rect 289078 158760 289084 158772
rect 160980 158732 289084 158760
rect 160980 158720 160986 158732
rect 289078 158720 289084 158732
rect 289136 158720 289142 158772
rect 297818 158720 297824 158772
rect 297876 158760 297882 158772
rect 373350 158760 373356 158772
rect 297876 158732 373356 158760
rect 297876 158720 297882 158732
rect 373350 158720 373356 158732
rect 373408 158720 373414 158772
rect 120626 158652 120632 158704
rect 120684 158692 120690 158704
rect 288066 158692 288072 158704
rect 120684 158664 288072 158692
rect 120684 158652 120690 158664
rect 288066 158652 288072 158664
rect 288124 158692 288130 158704
rect 288250 158692 288256 158704
rect 288124 158664 288256 158692
rect 288124 158652 288130 158664
rect 288250 158652 288256 158664
rect 288308 158652 288314 158704
rect 290826 158652 290832 158704
rect 290884 158692 290890 158704
rect 340966 158692 340972 158704
rect 290884 158664 340972 158692
rect 290884 158652 290890 158664
rect 340966 158652 340972 158664
rect 341024 158652 341030 158704
rect 376018 158652 376024 158704
rect 376076 158692 376082 158704
rect 438026 158692 438032 158704
rect 376076 158664 438032 158692
rect 376076 158652 376082 158664
rect 438026 158652 438032 158664
rect 438084 158652 438090 158704
rect 282546 158584 282552 158636
rect 282604 158624 282610 158636
rect 345934 158624 345940 158636
rect 282604 158596 345940 158624
rect 282604 158584 282610 158596
rect 345934 158584 345940 158596
rect 345992 158584 345998 158636
rect 378594 158584 378600 158636
rect 378652 158624 378658 158636
rect 439498 158624 439504 158636
rect 378652 158596 439504 158624
rect 378652 158584 378658 158596
rect 439498 158584 439504 158596
rect 439556 158584 439562 158636
rect 119706 158516 119712 158568
rect 119764 158556 119770 158568
rect 286134 158556 286140 158568
rect 119764 158528 286140 158556
rect 119764 158516 119770 158528
rect 286134 158516 286140 158528
rect 286192 158556 286198 158568
rect 286686 158556 286692 158568
rect 286192 158528 286692 158556
rect 286192 158516 286198 158528
rect 286686 158516 286692 158528
rect 286744 158516 286750 158568
rect 286778 158516 286784 158568
rect 286836 158556 286842 158568
rect 365806 158556 365812 158568
rect 286836 158528 365812 158556
rect 286836 158516 286842 158528
rect 365806 158516 365812 158528
rect 365864 158516 365870 158568
rect 380986 158516 380992 158568
rect 381044 158556 381050 158568
rect 436830 158556 436836 158568
rect 381044 158528 436836 158556
rect 381044 158516 381050 158528
rect 436830 158516 436836 158528
rect 436888 158516 436894 158568
rect 288158 158448 288164 158500
rect 288216 158488 288222 158500
rect 343542 158488 343548 158500
rect 288216 158460 343548 158488
rect 288216 158448 288222 158460
rect 343542 158448 343548 158460
rect 343600 158448 343606 158500
rect 383562 158448 383568 158500
rect 383620 158488 383626 158500
rect 438118 158488 438124 158500
rect 383620 158460 438124 158488
rect 383620 158448 383626 158460
rect 438118 158448 438124 158460
rect 438176 158448 438182 158500
rect 126514 158380 126520 158432
rect 126572 158420 126578 158432
rect 292298 158420 292304 158432
rect 126572 158392 292304 158420
rect 126572 158380 126578 158392
rect 292298 158380 292304 158392
rect 292356 158380 292362 158432
rect 293678 158380 293684 158432
rect 293736 158420 293742 158432
rect 328270 158420 328276 158432
rect 293736 158392 328276 158420
rect 293736 158380 293742 158392
rect 328270 158380 328276 158392
rect 328328 158380 328334 158432
rect 385954 158380 385960 158432
rect 386012 158420 386018 158432
rect 439590 158420 439596 158432
rect 386012 158392 439596 158420
rect 386012 158380 386018 158392
rect 439590 158380 439596 158392
rect 439648 158380 439654 158432
rect 133506 158312 133512 158364
rect 133564 158352 133570 158364
rect 299198 158352 299204 158364
rect 133564 158324 299204 158352
rect 133564 158312 133570 158324
rect 299198 158312 299204 158324
rect 299256 158352 299262 158364
rect 333422 158352 333428 158364
rect 299256 158324 333428 158352
rect 299256 158312 299262 158324
rect 333422 158312 333428 158324
rect 333480 158312 333486 158364
rect 388530 158312 388536 158364
rect 388588 158352 388594 158364
rect 436922 158352 436928 158364
rect 388588 158324 436928 158352
rect 388588 158312 388594 158324
rect 436922 158312 436928 158324
rect 436980 158312 436986 158364
rect 130562 158244 130568 158296
rect 130620 158284 130626 158296
rect 281442 158284 281448 158296
rect 130620 158256 281448 158284
rect 130620 158244 130626 158256
rect 281442 158244 281448 158256
rect 281500 158284 281506 158296
rect 329926 158284 329932 158296
rect 281500 158256 329932 158284
rect 281500 158244 281506 158256
rect 329926 158244 329932 158256
rect 329984 158244 329990 158296
rect 391474 158244 391480 158296
rect 391532 158284 391538 158296
rect 438302 158284 438308 158296
rect 391532 158256 438308 158284
rect 391532 158244 391538 158256
rect 438302 158244 438308 158256
rect 438360 158244 438366 158296
rect 128170 158176 128176 158228
rect 128228 158216 128234 158228
rect 274358 158216 274364 158228
rect 128228 158188 274364 158216
rect 128228 158176 128234 158188
rect 274358 158176 274364 158188
rect 274416 158176 274422 158228
rect 285398 158176 285404 158228
rect 285456 158216 285462 158228
rect 330570 158216 330576 158228
rect 285456 158188 330576 158216
rect 285456 158176 285462 158188
rect 330570 158176 330576 158188
rect 330628 158176 330634 158228
rect 394234 158176 394240 158228
rect 394292 158216 394298 158228
rect 440602 158216 440608 158228
rect 394292 158188 440608 158216
rect 394292 158176 394298 158188
rect 440602 158176 440608 158188
rect 440660 158176 440666 158228
rect 128722 158108 128728 158160
rect 128780 158148 128786 158160
rect 274450 158148 274456 158160
rect 128780 158120 274456 158148
rect 128780 158108 128786 158120
rect 274450 158108 274456 158120
rect 274508 158108 274514 158160
rect 292298 158108 292304 158160
rect 292356 158148 292362 158160
rect 326430 158148 326436 158160
rect 292356 158120 326436 158148
rect 292356 158108 292362 158120
rect 326430 158108 326436 158120
rect 326488 158108 326494 158160
rect 395890 158108 395896 158160
rect 395948 158148 395954 158160
rect 441890 158148 441896 158160
rect 395948 158120 441896 158148
rect 395948 158108 395954 158120
rect 441890 158108 441896 158120
rect 441948 158108 441954 158160
rect 131482 158040 131488 158092
rect 131540 158080 131546 158092
rect 271690 158080 271696 158092
rect 131540 158052 271696 158080
rect 131540 158040 131546 158052
rect 271690 158040 271696 158052
rect 271748 158040 271754 158092
rect 285490 158080 285496 158092
rect 283300 158052 285496 158080
rect 132402 157972 132408 158024
rect 132460 158012 132466 158024
rect 271598 158012 271604 158024
rect 132460 157984 271604 158012
rect 132460 157972 132466 157984
rect 271598 157972 271604 157984
rect 271656 157972 271662 158024
rect 158530 157904 158536 157956
rect 158588 157944 158594 157956
rect 276014 157944 276020 157956
rect 158588 157916 276020 157944
rect 158588 157904 158594 157916
rect 276014 157904 276020 157916
rect 276072 157904 276078 157956
rect 159910 157836 159916 157888
rect 159968 157876 159974 157888
rect 271322 157876 271328 157888
rect 159968 157848 271328 157876
rect 159968 157836 159974 157848
rect 271322 157836 271328 157848
rect 271380 157836 271386 157888
rect 271414 157836 271420 157888
rect 271472 157876 271478 157888
rect 277946 157876 277952 157888
rect 271472 157848 277952 157876
rect 271472 157836 271478 157848
rect 277946 157836 277952 157848
rect 278004 157836 278010 157888
rect 234614 157768 234620 157820
rect 234672 157808 234678 157820
rect 283300 157808 283328 158052
rect 285490 158040 285496 158052
rect 285548 158080 285554 158092
rect 318150 158080 318156 158092
rect 285548 158052 318156 158080
rect 285548 158040 285554 158052
rect 318150 158040 318156 158052
rect 318208 158040 318214 158092
rect 398466 158040 398472 158092
rect 398524 158080 398530 158092
rect 441798 158080 441804 158092
rect 398524 158052 441804 158080
rect 398524 158040 398530 158052
rect 441798 158040 441804 158052
rect 441856 158040 441862 158092
rect 289354 157972 289360 158024
rect 289412 158012 289418 158024
rect 289538 158012 289544 158024
rect 289412 157984 289544 158012
rect 289412 157972 289418 157984
rect 289538 157972 289544 157984
rect 289596 158012 289602 158024
rect 321646 158012 321652 158024
rect 289596 157984 321652 158012
rect 289596 157972 289602 157984
rect 321646 157972 321652 157984
rect 321704 157972 321710 158024
rect 401042 157972 401048 158024
rect 401100 158012 401106 158024
rect 441706 158012 441712 158024
rect 401100 157984 441712 158012
rect 401100 157972 401106 157984
rect 441706 157972 441712 157984
rect 441764 157972 441770 158024
rect 286134 157904 286140 157956
rect 286192 157944 286198 157956
rect 319438 157944 319444 157956
rect 286192 157916 319444 157944
rect 286192 157904 286198 157916
rect 319438 157904 319444 157916
rect 319496 157904 319502 157956
rect 403986 157904 403992 157956
rect 404044 157944 404050 157956
rect 438210 157944 438216 157956
rect 404044 157916 438216 157944
rect 404044 157904 404050 157916
rect 438210 157904 438216 157916
rect 438268 157904 438274 157956
rect 288250 157836 288256 157888
rect 288308 157876 288314 157888
rect 320542 157876 320548 157888
rect 288308 157848 320548 157876
rect 288308 157836 288314 157848
rect 320542 157836 320548 157848
rect 320600 157836 320606 157888
rect 406470 157836 406476 157888
rect 406528 157876 406534 157888
rect 439682 157876 439688 157888
rect 406528 157848 439688 157876
rect 406528 157836 406534 157848
rect 439682 157836 439688 157848
rect 439740 157836 439746 157888
rect 234672 157780 258074 157808
rect 234672 157768 234678 157780
rect 258046 157740 258074 157780
rect 271432 157780 283328 157808
rect 271432 157740 271460 157780
rect 258046 157712 271460 157740
rect 97626 157632 97632 157684
rect 97684 157672 97690 157684
rect 297358 157672 297364 157684
rect 97684 157644 297364 157672
rect 97684 157632 97690 157644
rect 297358 157632 297364 157644
rect 297416 157632 297422 157684
rect 121914 157564 121920 157616
rect 121972 157604 121978 157616
rect 289354 157604 289360 157616
rect 121972 157576 289360 157604
rect 121972 157564 121978 157576
rect 289354 157564 289360 157576
rect 289412 157564 289418 157616
rect 271322 157496 271328 157548
rect 271380 157536 271386 157548
rect 274634 157536 274640 157548
rect 271380 157508 274640 157536
rect 271380 157496 271386 157508
rect 274634 157496 274640 157508
rect 274692 157496 274698 157548
rect 329742 157428 329748 157480
rect 329800 157468 329806 157480
rect 355226 157468 355232 157480
rect 329800 157440 355232 157468
rect 329800 157428 329806 157440
rect 355226 157428 355232 157440
rect 355284 157428 355290 157480
rect 321554 157360 321560 157412
rect 321612 157400 321618 157412
rect 356974 157400 356980 157412
rect 321612 157372 356980 157400
rect 321612 157360 321618 157372
rect 356974 157360 356980 157372
rect 357032 157360 357038 157412
rect 123202 157292 123208 157344
rect 123260 157332 123266 157344
rect 290734 157332 290740 157344
rect 123260 157304 290740 157332
rect 123260 157292 123266 157304
rect 290734 157292 290740 157304
rect 290792 157292 290798 157344
rect 295702 157292 295708 157344
rect 295760 157332 295766 157344
rect 296346 157332 296352 157344
rect 295760 157304 296352 157332
rect 295760 157292 295766 157304
rect 296346 157292 296352 157304
rect 296404 157332 296410 157344
rect 343910 157332 343916 157344
rect 296404 157304 343916 157332
rect 296404 157292 296410 157304
rect 343910 157292 343916 157304
rect 343968 157292 343974 157344
rect 273714 157224 273720 157276
rect 273772 157264 273778 157276
rect 274174 157264 274180 157276
rect 273772 157236 274180 157264
rect 273772 157224 273778 157236
rect 274174 157224 274180 157236
rect 274232 157264 274238 157276
rect 348694 157264 348700 157276
rect 274232 157236 348700 157264
rect 274232 157224 274238 157236
rect 348694 157224 348700 157236
rect 348752 157224 348758 157276
rect 117314 157156 117320 157208
rect 117372 157196 117378 157208
rect 282730 157196 282736 157208
rect 117372 157168 282736 157196
rect 117372 157156 117378 157168
rect 282730 157156 282736 157168
rect 282788 157156 282794 157208
rect 286870 157156 286876 157208
rect 286928 157196 286934 157208
rect 333606 157196 333612 157208
rect 286928 157168 333612 157196
rect 286928 157156 286934 157168
rect 333606 157156 333612 157168
rect 333664 157156 333670 157208
rect 116486 157088 116492 157140
rect 116544 157128 116550 157140
rect 282822 157128 282828 157140
rect 116544 157100 282828 157128
rect 116544 157088 116550 157100
rect 282822 157088 282828 157100
rect 282880 157128 282886 157140
rect 316034 157128 316040 157140
rect 282880 157100 316040 157128
rect 282880 157088 282886 157100
rect 316034 157088 316040 157100
rect 316092 157088 316098 157140
rect 134886 157020 134892 157072
rect 134944 157060 134950 157072
rect 279970 157060 279976 157072
rect 134944 157032 279976 157060
rect 134944 157020 134950 157032
rect 279970 157020 279976 157032
rect 280028 157060 280034 157072
rect 334526 157060 334532 157072
rect 280028 157032 334532 157060
rect 280028 157020 280034 157032
rect 334526 157020 334532 157032
rect 334584 157020 334590 157072
rect 135898 156952 135904 157004
rect 135956 156992 135962 157004
rect 277210 156992 277216 157004
rect 135956 156964 277216 156992
rect 135956 156952 135962 156964
rect 277210 156952 277216 156964
rect 277268 156992 277274 157004
rect 335630 156992 335636 157004
rect 277268 156964 335636 156992
rect 277268 156952 277274 156964
rect 335630 156952 335636 156964
rect 335688 156952 335694 157004
rect 138106 156884 138112 156936
rect 138164 156924 138170 156936
rect 277118 156924 277124 156936
rect 138164 156896 277124 156924
rect 138164 156884 138170 156896
rect 277118 156884 277124 156896
rect 277176 156924 277182 156936
rect 338114 156924 338120 156936
rect 277176 156896 338120 156924
rect 277176 156884 277182 156896
rect 338114 156884 338120 156896
rect 338172 156884 338178 156936
rect 137002 156816 137008 156868
rect 137060 156856 137066 156868
rect 274542 156856 274548 156868
rect 137060 156828 274548 156856
rect 137060 156816 137066 156828
rect 274542 156816 274548 156828
rect 274600 156856 274606 156868
rect 336826 156856 336832 156868
rect 274600 156828 336832 156856
rect 274600 156816 274606 156828
rect 336826 156816 336832 156828
rect 336884 156816 336890 156868
rect 148870 156748 148876 156800
rect 148928 156788 148934 156800
rect 273714 156788 273720 156800
rect 148928 156760 273720 156788
rect 148928 156748 148934 156760
rect 273714 156748 273720 156760
rect 273772 156748 273778 156800
rect 282730 156748 282736 156800
rect 282788 156788 282794 156800
rect 316954 156788 316960 156800
rect 282788 156760 316960 156788
rect 282788 156748 282794 156760
rect 316954 156748 316960 156760
rect 317012 156748 317018 156800
rect 118234 156680 118240 156732
rect 118292 156720 118298 156732
rect 234614 156720 234620 156732
rect 118292 156692 234620 156720
rect 118292 156680 118298 156692
rect 234614 156680 234620 156692
rect 234672 156680 234678 156732
rect 287422 156680 287428 156732
rect 287480 156720 287486 156732
rect 306374 156720 306380 156732
rect 287480 156692 306380 156720
rect 287480 156680 287486 156692
rect 306374 156680 306380 156692
rect 306432 156680 306438 156732
rect 178862 156612 178868 156664
rect 178920 156652 178926 156664
rect 275370 156652 275376 156664
rect 178920 156624 275376 156652
rect 178920 156612 178926 156624
rect 275370 156612 275376 156624
rect 275428 156612 275434 156664
rect 291930 156612 291936 156664
rect 291988 156652 291994 156664
rect 313274 156652 313280 156664
rect 291988 156624 313280 156652
rect 291988 156612 291994 156624
rect 313274 156612 313280 156624
rect 313332 156612 313338 156664
rect 181806 156544 181812 156596
rect 181864 156584 181870 156596
rect 275278 156584 275284 156596
rect 181864 156556 275284 156584
rect 181864 156544 181870 156556
rect 275278 156544 275284 156556
rect 275336 156544 275342 156596
rect 290734 156544 290740 156596
rect 290792 156584 290798 156596
rect 323118 156584 323124 156596
rect 290792 156556 323124 156584
rect 290792 156544 290798 156556
rect 323118 156544 323124 156556
rect 323176 156544 323182 156596
rect 184014 156476 184020 156528
rect 184072 156516 184078 156528
rect 272518 156516 272524 156528
rect 184072 156488 272524 156516
rect 184072 156476 184078 156488
rect 272518 156476 272524 156488
rect 272576 156476 272582 156528
rect 185946 156408 185952 156460
rect 186004 156448 186010 156460
rect 272610 156448 272616 156460
rect 186004 156420 272616 156448
rect 186004 156408 186010 156420
rect 272610 156408 272616 156420
rect 272668 156408 272674 156460
rect 144086 156340 144092 156392
rect 144144 156380 144150 156392
rect 295702 156380 295708 156392
rect 144144 156352 295708 156380
rect 144144 156340 144150 156352
rect 295702 156340 295708 156352
rect 295760 156340 295766 156392
rect 280062 155864 280068 155916
rect 280120 155904 280126 155916
rect 338206 155904 338212 155916
rect 280120 155876 338212 155904
rect 280120 155864 280126 155876
rect 338206 155864 338212 155876
rect 338264 155864 338270 155916
rect 140682 155796 140688 155848
rect 140740 155836 140746 155848
rect 284110 155836 284116 155848
rect 140740 155808 284116 155836
rect 140740 155796 140746 155808
rect 284110 155796 284116 155808
rect 284168 155836 284174 155848
rect 339494 155836 339500 155848
rect 284168 155808 339500 155836
rect 284168 155796 284174 155808
rect 339494 155796 339500 155808
rect 339552 155796 339558 155848
rect 274634 155728 274640 155780
rect 274692 155768 274698 155780
rect 275830 155768 275836 155780
rect 274692 155740 275836 155768
rect 274692 155728 274698 155740
rect 275830 155728 275836 155740
rect 275888 155768 275894 155780
rect 346670 155768 346676 155780
rect 275888 155740 346676 155768
rect 275888 155728 275894 155740
rect 346670 155728 346676 155740
rect 346728 155728 346734 155780
rect 294322 155660 294328 155712
rect 294380 155700 294386 155712
rect 294966 155700 294972 155712
rect 294380 155672 294972 155700
rect 294380 155660 294386 155672
rect 294966 155660 294972 155672
rect 295024 155700 295030 155712
rect 342346 155700 342352 155712
rect 295024 155672 342352 155700
rect 295024 155660 295030 155672
rect 342346 155660 342352 155672
rect 342404 155660 342410 155712
rect 140498 155592 140504 155644
rect 140556 155632 140562 155644
rect 280062 155632 280068 155644
rect 140556 155604 280068 155632
rect 140556 155592 140562 155604
rect 280062 155592 280068 155604
rect 280120 155592 280126 155644
rect 281442 155592 281448 155644
rect 281500 155632 281506 155644
rect 345106 155632 345112 155644
rect 281500 155604 345112 155632
rect 281500 155592 281506 155604
rect 345106 155592 345112 155604
rect 345164 155592 345170 155644
rect 141786 155524 141792 155576
rect 141844 155564 141850 155576
rect 278590 155564 278596 155576
rect 141844 155536 278596 155564
rect 141844 155524 141850 155536
rect 278590 155524 278596 155536
rect 278648 155564 278654 155576
rect 341058 155564 341064 155576
rect 278648 155536 341064 155564
rect 278648 155524 278654 155536
rect 341058 155524 341064 155536
rect 341116 155524 341122 155576
rect 145282 155456 145288 155508
rect 145340 155496 145346 155508
rect 281442 155496 281448 155508
rect 145340 155468 281448 155496
rect 145340 155456 145346 155468
rect 281442 155456 281448 155468
rect 281500 155456 281506 155508
rect 295702 155456 295708 155508
rect 295760 155496 295766 155508
rect 296530 155496 296536 155508
rect 295760 155468 296536 155496
rect 295760 155456 295766 155468
rect 296530 155456 296536 155468
rect 296588 155496 296594 155508
rect 324222 155496 324228 155508
rect 296588 155468 324228 155496
rect 296588 155456 296594 155468
rect 324222 155456 324228 155468
rect 324280 155456 324286 155508
rect 146386 155388 146392 155440
rect 146444 155428 146450 155440
rect 277302 155428 277308 155440
rect 146444 155400 277308 155428
rect 146444 155388 146450 155400
rect 277302 155388 277308 155400
rect 277360 155428 277366 155440
rect 346394 155428 346400 155440
rect 277360 155400 346400 155428
rect 277360 155388 277366 155400
rect 346394 155388 346400 155400
rect 346452 155388 346458 155440
rect 136082 155320 136088 155372
rect 136140 155360 136146 155372
rect 265710 155360 265716 155372
rect 136140 155332 265716 155360
rect 136140 155320 136146 155332
rect 265710 155320 265716 155332
rect 265768 155320 265774 155372
rect 299290 155320 299296 155372
rect 299348 155360 299354 155372
rect 321554 155360 321560 155372
rect 299348 155332 321560 155360
rect 299348 155320 299354 155332
rect 321554 155320 321560 155332
rect 321612 155320 321618 155372
rect 147674 155252 147680 155304
rect 147732 155292 147738 155304
rect 274634 155292 274640 155304
rect 147732 155264 274640 155292
rect 147732 155252 147738 155264
rect 274634 155252 274640 155264
rect 274692 155252 274698 155304
rect 195882 155184 195888 155236
rect 195940 155224 195946 155236
rect 266998 155224 267004 155236
rect 195940 155196 267004 155224
rect 195940 155184 195946 155196
rect 266998 155184 267004 155196
rect 267056 155184 267062 155236
rect 198458 155116 198464 155168
rect 198516 155156 198522 155168
rect 267182 155156 267188 155168
rect 198516 155128 267188 155156
rect 198516 155116 198522 155128
rect 267182 155116 267188 155128
rect 267240 155116 267246 155168
rect 201034 155048 201040 155100
rect 201092 155088 201098 155100
rect 264330 155088 264336 155100
rect 201092 155060 264336 155088
rect 201092 155048 201098 155060
rect 264330 155048 264336 155060
rect 264388 155048 264394 155100
rect 203426 154980 203432 155032
rect 203484 155020 203490 155032
rect 261570 155020 261576 155032
rect 203484 154992 261576 155020
rect 203484 154980 203490 154992
rect 261570 154980 261576 154992
rect 261628 154980 261634 155032
rect 124582 154912 124588 154964
rect 124640 154952 124646 154964
rect 295702 154952 295708 154964
rect 124640 154924 295708 154952
rect 124640 154912 124646 154924
rect 295702 154912 295708 154924
rect 295760 154912 295766 154964
rect 143074 154844 143080 154896
rect 143132 154884 143138 154896
rect 294322 154884 294328 154896
rect 143132 154856 294328 154884
rect 143132 154844 143138 154856
rect 294322 154844 294328 154856
rect 294380 154844 294386 154896
rect 157058 154776 157064 154828
rect 157116 154816 157122 154828
rect 298370 154816 298376 154828
rect 157116 154788 298376 154816
rect 157116 154776 157122 154788
rect 298370 154776 298376 154788
rect 298428 154816 298434 154828
rect 299290 154816 299296 154828
rect 298428 154788 299296 154816
rect 298428 154776 298434 154788
rect 299290 154776 299296 154788
rect 299348 154776 299354 154828
rect 284754 154572 284760 154624
rect 284812 154612 284818 154624
rect 287422 154612 287428 154624
rect 284812 154584 287428 154612
rect 284812 154572 284818 154584
rect 287422 154572 287428 154584
rect 287480 154572 287486 154624
rect 125410 154504 125416 154556
rect 125468 154544 125474 154556
rect 271782 154544 271788 154556
rect 125468 154516 271788 154544
rect 125468 154504 125474 154516
rect 271782 154504 271788 154516
rect 271840 154504 271846 154556
rect 272702 154504 272708 154556
rect 272760 154544 272766 154556
rect 273162 154544 273168 154556
rect 272760 154516 273168 154544
rect 272760 154504 272766 154516
rect 273162 154504 273168 154516
rect 273220 154544 273226 154556
rect 354398 154544 354404 154556
rect 273220 154516 354404 154544
rect 273220 154504 273226 154516
rect 354398 154504 354404 154516
rect 354456 154504 354462 154556
rect 154114 154436 154120 154488
rect 154172 154476 154178 154488
rect 298002 154476 298008 154488
rect 154172 154448 298008 154476
rect 154172 154436 154178 154448
rect 298002 154436 298008 154448
rect 298060 154476 298066 154488
rect 353294 154476 353300 154488
rect 298060 154448 353300 154476
rect 298060 154436 298066 154448
rect 353294 154436 353300 154448
rect 353352 154436 353358 154488
rect 155770 154368 155776 154420
rect 155828 154408 155834 154420
rect 298554 154408 298560 154420
rect 155828 154380 298560 154408
rect 155828 154368 155834 154380
rect 298554 154368 298560 154380
rect 298612 154408 298618 154420
rect 329742 154408 329748 154420
rect 298612 154380 329748 154408
rect 298612 154368 298618 154380
rect 329742 154368 329748 154380
rect 329800 154368 329806 154420
rect 152642 154300 152648 154352
rect 152700 154340 152706 154352
rect 284202 154340 284208 154352
rect 152700 154312 284208 154340
rect 152700 154300 152706 154312
rect 284202 154300 284208 154312
rect 284260 154340 284266 154352
rect 352190 154340 352196 154352
rect 284260 154312 352196 154340
rect 284260 154300 284266 154312
rect 352190 154300 352196 154312
rect 352248 154300 352254 154352
rect 149882 154232 149888 154284
rect 149940 154272 149946 154284
rect 279878 154272 279884 154284
rect 149940 154244 279884 154272
rect 149940 154232 149946 154244
rect 279878 154232 279884 154244
rect 279936 154272 279942 154284
rect 349798 154272 349804 154284
rect 279936 154244 349804 154272
rect 279936 154232 279942 154244
rect 349798 154232 349804 154244
rect 349856 154232 349862 154284
rect 151354 154164 151360 154216
rect 151412 154204 151418 154216
rect 278682 154204 278688 154216
rect 151412 154176 278688 154204
rect 151412 154164 151418 154176
rect 278682 154164 278688 154176
rect 278740 154204 278746 154216
rect 350994 154204 351000 154216
rect 278740 154176 351000 154204
rect 278740 154164 278746 154176
rect 350994 154164 351000 154176
rect 351052 154164 351058 154216
rect 271782 154096 271788 154148
rect 271840 154136 271846 154148
rect 325326 154136 325332 154148
rect 271840 154108 325332 154136
rect 271840 154096 271846 154108
rect 325326 154096 325332 154108
rect 325384 154096 325390 154148
rect 227714 154028 227720 154080
rect 227772 154068 227778 154080
rect 275002 154068 275008 154080
rect 227772 154040 275008 154068
rect 227772 154028 227778 154040
rect 275002 154028 275008 154040
rect 275060 154028 275066 154080
rect 208394 153960 208400 154012
rect 208452 154000 208458 154012
rect 272334 154000 272340 154012
rect 208452 153972 272340 154000
rect 208452 153960 208458 153972
rect 272334 153960 272340 153972
rect 272392 153960 272398 154012
rect 193214 153892 193220 153944
rect 193272 153932 193278 153944
rect 269666 153932 269672 153944
rect 193272 153904 269672 153932
rect 193272 153892 193278 153904
rect 269666 153892 269672 153904
rect 269724 153892 269730 153944
rect 286042 153892 286048 153944
rect 286100 153932 286106 153944
rect 292942 153932 292948 153944
rect 286100 153904 292948 153932
rect 286100 153892 286106 153904
rect 292942 153892 292948 153904
rect 293000 153892 293006 153944
rect 168374 153824 168380 153876
rect 168432 153864 168438 153876
rect 265434 153864 265440 153876
rect 168432 153836 265440 153864
rect 168432 153824 168438 153836
rect 265434 153824 265440 153836
rect 265492 153824 265498 153876
rect 287330 153824 287336 153876
rect 287388 153864 287394 153876
rect 304994 153864 305000 153876
rect 287388 153836 305000 153864
rect 287388 153824 287394 153836
rect 304994 153824 305000 153836
rect 305052 153824 305058 153876
rect 154482 153756 154488 153808
rect 154540 153796 154546 153808
rect 272702 153796 272708 153808
rect 154540 153768 272708 153796
rect 154540 153756 154546 153768
rect 272702 153756 272708 153768
rect 272760 153756 272766 153808
rect 141418 153144 141424 153196
rect 141476 153184 141482 153196
rect 258902 153184 258908 153196
rect 141476 153156 258908 153184
rect 141476 153144 141482 153156
rect 258902 153144 258908 153156
rect 258960 153144 258966 153196
rect 144362 153076 144368 153128
rect 144420 153116 144426 153128
rect 258810 153116 258816 153128
rect 144420 153088 258816 153116
rect 144420 153076 144426 153088
rect 258810 153076 258816 153088
rect 258868 153076 258874 153128
rect 146018 153008 146024 153060
rect 146076 153048 146082 153060
rect 258718 153048 258724 153060
rect 146076 153020 258724 153048
rect 146076 153008 146082 153020
rect 258718 153008 258724 153020
rect 258776 153008 258782 153060
rect 148502 152940 148508 152992
rect 148560 152980 148566 152992
rect 256142 152980 256148 152992
rect 148560 152952 256148 152980
rect 148560 152940 148566 152952
rect 256142 152940 256148 152952
rect 256200 152940 256206 152992
rect 150986 152872 150992 152924
rect 151044 152912 151050 152924
rect 256234 152912 256240 152924
rect 151044 152884 256240 152912
rect 151044 152872 151050 152884
rect 256234 152872 256240 152884
rect 256292 152872 256298 152924
rect 288894 152668 288900 152720
rect 288952 152708 288958 152720
rect 310514 152708 310520 152720
rect 288952 152680 310520 152708
rect 288952 152668 288958 152680
rect 310514 152668 310520 152680
rect 310572 152668 310578 152720
rect 291654 152600 291660 152652
rect 291712 152640 291718 152652
rect 331214 152640 331220 152652
rect 291712 152612 331220 152640
rect 291712 152600 291718 152612
rect 331214 152600 331220 152612
rect 331272 152600 331278 152652
rect 295610 152532 295616 152584
rect 295668 152572 295674 152584
rect 357434 152572 357440 152584
rect 295668 152544 357440 152572
rect 295668 152532 295674 152544
rect 357434 152532 357440 152544
rect 357492 152532 357498 152584
rect 135254 152464 135260 152516
rect 135312 152504 135318 152516
rect 261478 152504 261484 152516
rect 135312 152476 261484 152504
rect 135312 152464 135318 152476
rect 261478 152464 261484 152476
rect 261536 152464 261542 152516
rect 271230 152464 271236 152516
rect 271288 152504 271294 152516
rect 280430 152504 280436 152516
rect 271288 152476 280436 152504
rect 271288 152464 271294 152476
rect 280430 152464 280436 152476
rect 280488 152464 280494 152516
rect 298186 152464 298192 152516
rect 298244 152504 298250 152516
rect 374086 152504 374092 152516
rect 298244 152476 374092 152504
rect 298244 152464 298250 152476
rect 374086 152464 374092 152476
rect 374144 152464 374150 152516
rect 182174 151104 182180 151156
rect 182232 151144 182238 151156
rect 268194 151144 268200 151156
rect 182232 151116 268200 151144
rect 182232 151104 182238 151116
rect 268194 151104 268200 151116
rect 268252 151104 268258 151156
rect 285950 151104 285956 151156
rect 286008 151144 286014 151156
rect 299566 151144 299572 151156
rect 286008 151116 299572 151144
rect 286008 151104 286014 151116
rect 299566 151104 299572 151116
rect 299624 151104 299630 151156
rect 146294 151036 146300 151088
rect 146352 151076 146358 151088
rect 262582 151076 262588 151088
rect 146352 151048 262588 151076
rect 146352 151036 146358 151048
rect 262582 151036 262588 151048
rect 262640 151036 262646 151088
rect 291562 151036 291568 151088
rect 291620 151076 291626 151088
rect 333974 151076 333980 151088
rect 291620 151048 333980 151076
rect 291620 151036 291626 151048
rect 333974 151036 333980 151048
rect 334032 151036 334038 151088
rect 184934 149812 184940 149864
rect 184992 149852 184998 149864
rect 268102 149852 268108 149864
rect 184992 149824 268108 149852
rect 184992 149812 184998 149824
rect 268102 149812 268108 149824
rect 268160 149812 268166 149864
rect 157334 149744 157340 149796
rect 157392 149784 157398 149796
rect 264146 149784 264152 149796
rect 157392 149756 264152 149784
rect 157392 149744 157398 149756
rect 264146 149744 264152 149756
rect 264204 149744 264210 149796
rect 288802 149744 288808 149796
rect 288860 149784 288866 149796
rect 314654 149784 314660 149796
rect 288860 149756 314660 149784
rect 288860 149744 288866 149756
rect 314654 149744 314660 149756
rect 314712 149744 314718 149796
rect 121454 149676 121460 149728
rect 121512 149716 121518 149728
rect 258442 149716 258448 149728
rect 121512 149688 258448 149716
rect 121512 149676 121518 149688
rect 258442 149676 258448 149688
rect 258500 149676 258506 149728
rect 292850 149676 292856 149728
rect 292908 149716 292914 149728
rect 340874 149716 340880 149728
rect 292908 149688 340880 149716
rect 292908 149676 292914 149688
rect 340874 149676 340880 149688
rect 340932 149676 340938 149728
rect 224954 148384 224960 148436
rect 225012 148424 225018 148436
rect 273898 148424 273904 148436
rect 225012 148396 273904 148424
rect 225012 148384 225018 148396
rect 273898 148384 273904 148396
rect 273956 148384 273962 148436
rect 128354 148316 128360 148368
rect 128412 148356 128418 148368
rect 259914 148356 259920 148368
rect 128412 148328 259920 148356
rect 128412 148316 128418 148328
rect 259914 148316 259920 148328
rect 259972 148316 259978 148368
rect 273990 148316 273996 148368
rect 274048 148356 274054 148368
rect 281994 148356 282000 148368
rect 274048 148328 282000 148356
rect 274048 148316 274054 148328
rect 281994 148316 282000 148328
rect 282052 148316 282058 148368
rect 285858 148316 285864 148368
rect 285916 148356 285922 148368
rect 300854 148356 300860 148368
rect 285916 148328 300860 148356
rect 285916 148316 285922 148328
rect 300854 148316 300860 148328
rect 300912 148316 300918 148368
rect 200114 146956 200120 147008
rect 200172 146996 200178 147008
rect 270862 146996 270868 147008
rect 200172 146968 270868 146996
rect 200172 146956 200178 146968
rect 270862 146956 270868 146968
rect 270920 146956 270926 147008
rect 281994 146956 282000 147008
rect 282052 146996 282058 147008
rect 283374 146996 283380 147008
rect 282052 146968 283380 146996
rect 282052 146956 282058 146968
rect 283374 146956 283380 146968
rect 283432 146956 283438 147008
rect 139394 146888 139400 146940
rect 139452 146928 139458 146940
rect 261386 146928 261392 146940
rect 139452 146900 261392 146928
rect 139452 146888 139458 146900
rect 261386 146888 261392 146900
rect 261444 146888 261450 146940
rect 270954 146888 270960 146940
rect 271012 146928 271018 146940
rect 281902 146928 281908 146940
rect 271012 146900 281908 146928
rect 271012 146888 271018 146900
rect 281902 146888 281908 146900
rect 281960 146888 281966 146940
rect 287238 146888 287244 146940
rect 287296 146928 287302 146940
rect 303614 146928 303620 146940
rect 287296 146900 303620 146928
rect 287296 146888 287302 146900
rect 303614 146888 303620 146900
rect 303672 146888 303678 146940
rect 218054 145664 218060 145716
rect 218112 145704 218118 145716
rect 273530 145704 273536 145716
rect 218112 145676 273536 145704
rect 218112 145664 218118 145676
rect 273530 145664 273536 145676
rect 273588 145664 273594 145716
rect 150434 145596 150440 145648
rect 150492 145636 150498 145648
rect 262490 145636 262496 145648
rect 150492 145608 262496 145636
rect 150492 145596 150498 145608
rect 262490 145596 262496 145608
rect 262548 145596 262554 145648
rect 133874 145528 133880 145580
rect 133932 145568 133938 145580
rect 261294 145568 261300 145580
rect 133932 145540 261300 145568
rect 133932 145528 133938 145540
rect 261294 145528 261300 145540
rect 261352 145528 261358 145580
rect 273898 145528 273904 145580
rect 273956 145568 273962 145580
rect 280338 145568 280344 145580
rect 273956 145540 280344 145568
rect 273956 145528 273962 145540
rect 280338 145528 280344 145540
rect 280396 145528 280402 145580
rect 288710 145528 288716 145580
rect 288768 145568 288774 145580
rect 317414 145568 317420 145580
rect 288768 145540 317420 145568
rect 288768 145528 288774 145540
rect 317414 145528 317420 145540
rect 317472 145528 317478 145580
rect 216674 144304 216680 144356
rect 216732 144344 216738 144356
rect 273438 144344 273444 144356
rect 216732 144316 273444 144344
rect 216732 144304 216738 144316
rect 273438 144304 273444 144316
rect 273496 144304 273502 144356
rect 186314 144236 186320 144288
rect 186372 144276 186378 144288
rect 269574 144276 269580 144288
rect 186372 144248 269580 144276
rect 186372 144236 186378 144248
rect 269574 144236 269580 144248
rect 269632 144236 269638 144288
rect 132494 144168 132500 144220
rect 132552 144208 132558 144220
rect 259822 144208 259828 144220
rect 132552 144180 259828 144208
rect 132552 144168 132558 144180
rect 259822 144168 259828 144180
rect 259880 144168 259886 144220
rect 260190 144168 260196 144220
rect 260248 144208 260254 144220
rect 279142 144208 279148 144220
rect 260248 144180 279148 144208
rect 260248 144168 260254 144180
rect 279142 144168 279148 144180
rect 279200 144168 279206 144220
rect 291470 144168 291476 144220
rect 291528 144208 291534 144220
rect 328454 144208 328460 144220
rect 291528 144180 328460 144208
rect 291528 144168 291534 144180
rect 328454 144168 328460 144180
rect 328512 144168 328518 144220
rect 209774 142944 209780 142996
rect 209832 142984 209838 142996
rect 272242 142984 272248 142996
rect 209832 142956 272248 142984
rect 209832 142944 209838 142956
rect 272242 142944 272248 142956
rect 272300 142944 272306 142996
rect 197354 142876 197360 142928
rect 197412 142916 197418 142928
rect 270770 142916 270776 142928
rect 197412 142888 270776 142916
rect 197412 142876 197418 142888
rect 270770 142876 270776 142888
rect 270828 142876 270834 142928
rect 286318 142876 286324 142928
rect 286376 142916 286382 142928
rect 291470 142916 291476 142928
rect 286376 142888 291476 142916
rect 286376 142876 286382 142888
rect 291470 142876 291476 142888
rect 291528 142876 291534 142928
rect 143534 142808 143540 142860
rect 143592 142848 143598 142860
rect 260098 142848 260104 142860
rect 143592 142820 260104 142848
rect 143592 142808 143598 142820
rect 260098 142808 260104 142820
rect 260156 142808 260162 142860
rect 291378 142808 291384 142860
rect 291436 142848 291442 142860
rect 332594 142848 332600 142860
rect 291436 142820 332600 142848
rect 291436 142808 291442 142820
rect 332594 142808 332600 142820
rect 332652 142808 332658 142860
rect 201494 141516 201500 141568
rect 201552 141556 201558 141568
rect 270678 141556 270684 141568
rect 201552 141528 270684 141556
rect 201552 141516 201558 141528
rect 270678 141516 270684 141528
rect 270736 141516 270742 141568
rect 126974 141448 126980 141500
rect 127032 141488 127038 141500
rect 259730 141488 259736 141500
rect 127032 141460 259736 141488
rect 127032 141448 127038 141460
rect 259730 141448 259736 141460
rect 259788 141448 259794 141500
rect 115934 141380 115940 141432
rect 115992 141420 115998 141432
rect 258350 141420 258356 141432
rect 115992 141392 258356 141420
rect 115992 141380 115998 141392
rect 258350 141380 258356 141392
rect 258408 141380 258414 141432
rect 291286 141380 291292 141432
rect 291344 141420 291350 141432
rect 335354 141420 335360 141432
rect 291344 141392 335360 141420
rect 291344 141380 291350 141392
rect 335354 141380 335360 141392
rect 335412 141380 335418 141432
rect 211154 140156 211160 140208
rect 211212 140196 211218 140208
rect 272150 140196 272156 140208
rect 211212 140168 272156 140196
rect 211212 140156 211218 140168
rect 272150 140156 272156 140168
rect 272208 140156 272214 140208
rect 161474 140088 161480 140140
rect 161532 140128 161538 140140
rect 265342 140128 265348 140140
rect 161532 140100 265348 140128
rect 161532 140088 161538 140100
rect 265342 140088 265348 140100
rect 265400 140088 265406 140140
rect 107654 140020 107660 140072
rect 107712 140060 107718 140072
rect 257062 140060 257068 140072
rect 107712 140032 257068 140060
rect 107712 140020 107718 140032
rect 257062 140020 257068 140032
rect 257120 140020 257126 140072
rect 292758 140020 292764 140072
rect 292816 140060 292822 140072
rect 339494 140060 339500 140072
rect 292816 140032 339500 140060
rect 292816 140020 292822 140032
rect 339494 140020 339500 140032
rect 339552 140020 339558 140072
rect 165614 138728 165620 138780
rect 165672 138768 165678 138780
rect 265250 138768 265256 138780
rect 165672 138740 265256 138768
rect 165672 138728 165678 138740
rect 265250 138728 265256 138740
rect 265308 138728 265314 138780
rect 110414 138660 110420 138712
rect 110472 138700 110478 138712
rect 256970 138700 256976 138712
rect 110472 138672 256976 138700
rect 110472 138660 110478 138672
rect 256970 138660 256976 138672
rect 257028 138660 257034 138712
rect 274082 138660 274088 138712
rect 274140 138700 274146 138712
rect 281810 138700 281816 138712
rect 274140 138672 281816 138700
rect 274140 138660 274146 138672
rect 281810 138660 281816 138672
rect 281868 138660 281874 138712
rect 292666 138660 292672 138712
rect 292724 138700 292730 138712
rect 342254 138700 342260 138712
rect 292724 138672 342260 138700
rect 292724 138660 292730 138672
rect 342254 138660 342260 138672
rect 342312 138660 342318 138712
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 84838 137952 84844 137964
rect 3568 137924 84844 137952
rect 3568 137912 3574 137924
rect 84838 137912 84844 137924
rect 84896 137912 84902 137964
rect 226334 137300 226340 137352
rect 226392 137340 226398 137352
rect 274910 137340 274916 137352
rect 226392 137312 274916 137340
rect 226392 137300 226398 137312
rect 274910 137300 274916 137312
rect 274968 137300 274974 137352
rect 103514 137232 103520 137284
rect 103572 137272 103578 137284
rect 255682 137272 255688 137284
rect 103572 137244 255688 137272
rect 103572 137232 103578 137244
rect 255682 137232 255688 137244
rect 255740 137232 255746 137284
rect 155954 135872 155960 135924
rect 156012 135912 156018 135924
rect 264054 135912 264060 135924
rect 156012 135884 264060 135912
rect 156012 135872 156018 135884
rect 264054 135872 264060 135884
rect 264112 135872 264118 135924
rect 179414 134580 179420 134632
rect 179472 134620 179478 134632
rect 268010 134620 268016 134632
rect 179472 134592 268016 134620
rect 179472 134580 179478 134592
rect 268010 134580 268016 134592
rect 268068 134580 268074 134632
rect 143626 134512 143632 134564
rect 143684 134552 143690 134564
rect 262398 134552 262404 134564
rect 143684 134524 262404 134552
rect 143684 134512 143690 134524
rect 262398 134512 262404 134524
rect 262456 134512 262462 134564
rect 266998 134512 267004 134564
rect 267056 134552 267062 134564
rect 280706 134552 280712 134564
rect 267056 134524 280712 134552
rect 267056 134512 267062 134524
rect 280706 134512 280712 134524
rect 280764 134512 280770 134564
rect 287146 134512 287152 134564
rect 287204 134552 287210 134564
rect 307754 134552 307760 134564
rect 287204 134524 307760 134552
rect 287204 134512 287210 134524
rect 307754 134512 307760 134524
rect 307812 134512 307818 134564
rect 183554 133220 183560 133272
rect 183612 133260 183618 133272
rect 267918 133260 267924 133272
rect 183612 133232 267924 133260
rect 183612 133220 183618 133232
rect 267918 133220 267924 133232
rect 267976 133220 267982 133272
rect 151814 133152 151820 133204
rect 151872 133192 151878 133204
rect 263962 133192 263968 133204
rect 151872 133164 263968 133192
rect 151872 133152 151878 133164
rect 263962 133152 263968 133164
rect 264020 133152 264026 133204
rect 268562 133152 268568 133204
rect 268620 133192 268626 133204
rect 279050 133192 279056 133204
rect 268620 133164 279056 133192
rect 268620 133152 268626 133164
rect 279050 133152 279056 133164
rect 279108 133152 279114 133204
rect 288618 133152 288624 133204
rect 288676 133192 288682 133204
rect 318794 133192 318800 133204
rect 288676 133164 318800 133192
rect 288676 133152 288682 133164
rect 318794 133152 318800 133164
rect 318852 133152 318858 133204
rect 187694 131792 187700 131844
rect 187752 131832 187758 131844
rect 265618 131832 265624 131844
rect 187752 131804 265624 131832
rect 187752 131792 187758 131804
rect 265618 131792 265624 131804
rect 265676 131792 265682 131844
rect 190454 131724 190460 131776
rect 190512 131764 190518 131776
rect 269482 131764 269488 131776
rect 190512 131736 269488 131764
rect 190512 131724 190518 131736
rect 269482 131724 269488 131736
rect 269540 131724 269546 131776
rect 293310 131724 293316 131776
rect 293368 131764 293374 131776
rect 332686 131764 332692 131776
rect 293368 131736 332692 131764
rect 293368 131724 293374 131736
rect 332686 131724 332692 131736
rect 332744 131724 332750 131776
rect 205634 130500 205640 130552
rect 205692 130540 205698 130552
rect 272058 130540 272064 130552
rect 205692 130512 272064 130540
rect 205692 130500 205698 130512
rect 272058 130500 272064 130512
rect 272116 130500 272122 130552
rect 193306 130432 193312 130484
rect 193364 130472 193370 130484
rect 269390 130472 269396 130484
rect 193364 130444 269396 130472
rect 193364 130432 193370 130444
rect 269390 130432 269396 130444
rect 269448 130432 269454 130484
rect 120074 130364 120080 130416
rect 120132 130404 120138 130416
rect 258258 130404 258264 130416
rect 120132 130376 258264 130404
rect 120132 130364 120138 130376
rect 258258 130364 258264 130376
rect 258316 130364 258322 130416
rect 292574 130364 292580 130416
rect 292632 130404 292638 130416
rect 340966 130404 340972 130416
rect 292632 130376 340972 130404
rect 292632 130364 292638 130376
rect 340966 130364 340972 130376
rect 341024 130364 341030 130416
rect 198734 129072 198740 129124
rect 198792 129112 198798 129124
rect 270586 129112 270592 129124
rect 198792 129084 270592 129112
rect 198792 129072 198798 129084
rect 270586 129072 270592 129084
rect 270644 129072 270650 129124
rect 129734 129004 129740 129056
rect 129792 129044 129798 129056
rect 259638 129044 259644 129056
rect 129792 129016 259644 129044
rect 129792 129004 129798 129016
rect 259638 129004 259644 129016
rect 259696 129004 259702 129056
rect 296162 129004 296168 129056
rect 296220 129044 296226 129056
rect 350534 129044 350540 129056
rect 296220 129016 350540 129044
rect 296220 129004 296226 129016
rect 350534 129004 350540 129016
rect 350592 129004 350598 129056
rect 204254 127644 204260 127696
rect 204312 127684 204318 127696
rect 271138 127684 271144 127696
rect 204312 127656 271144 127684
rect 204312 127644 204318 127656
rect 271138 127644 271144 127656
rect 271196 127644 271202 127696
rect 118694 127576 118700 127628
rect 118752 127616 118758 127628
rect 254578 127616 254584 127628
rect 118752 127588 254584 127616
rect 118752 127576 118758 127588
rect 254578 127576 254584 127588
rect 254636 127576 254642 127628
rect 218146 126284 218152 126336
rect 218204 126324 218210 126336
rect 273346 126324 273352 126336
rect 218204 126296 273352 126324
rect 218204 126284 218210 126296
rect 273346 126284 273352 126296
rect 273404 126284 273410 126336
rect 180794 126216 180800 126268
rect 180852 126256 180858 126268
rect 267826 126256 267832 126268
rect 180852 126228 267832 126256
rect 180852 126216 180858 126228
rect 267826 126216 267832 126228
rect 267884 126216 267890 126268
rect 229094 124924 229100 124976
rect 229152 124964 229158 124976
rect 274818 124964 274824 124976
rect 229152 124936 274824 124964
rect 229152 124924 229158 124936
rect 274818 124924 274824 124936
rect 274876 124924 274882 124976
rect 169754 124856 169760 124908
rect 169812 124896 169818 124908
rect 266722 124896 266728 124908
rect 169812 124868 266728 124896
rect 169812 124856 169818 124868
rect 266722 124856 266728 124868
rect 266780 124856 266786 124908
rect 275278 124856 275284 124908
rect 275336 124896 275342 124908
rect 281718 124896 281724 124908
rect 275336 124868 281724 124896
rect 275336 124856 275342 124868
rect 281718 124856 281724 124868
rect 281776 124856 281782 124908
rect 136634 123428 136640 123480
rect 136692 123468 136698 123480
rect 261202 123468 261208 123480
rect 136692 123440 261208 123468
rect 136692 123428 136698 123440
rect 261202 123428 261208 123440
rect 261260 123428 261266 123480
rect 140774 122068 140780 122120
rect 140832 122108 140838 122120
rect 261110 122108 261116 122120
rect 140832 122080 261116 122108
rect 140832 122068 140838 122080
rect 261110 122068 261116 122080
rect 261168 122068 261174 122120
rect 147674 120708 147680 120760
rect 147732 120748 147738 120760
rect 262306 120748 262312 120760
rect 147732 120720 262312 120748
rect 147732 120708 147738 120720
rect 262306 120708 262312 120720
rect 262364 120708 262370 120760
rect 154574 119348 154580 119400
rect 154632 119388 154638 119400
rect 263870 119388 263876 119400
rect 154632 119360 263876 119388
rect 154632 119348 154638 119360
rect 263870 119348 263876 119360
rect 263928 119348 263934 119400
rect 158714 117920 158720 117972
rect 158772 117960 158778 117972
rect 263778 117960 263784 117972
rect 158772 117932 263784 117960
rect 158772 117920 158778 117932
rect 263778 117920 263784 117932
rect 263836 117920 263842 117972
rect 127066 116560 127072 116612
rect 127124 116600 127130 116612
rect 259546 116600 259552 116612
rect 127124 116572 259552 116600
rect 127124 116560 127130 116572
rect 259546 116560 259552 116572
rect 259604 116560 259610 116612
rect 162854 115200 162860 115252
rect 162912 115240 162918 115252
rect 265158 115240 265164 115252
rect 162912 115212 265164 115240
rect 162912 115200 162918 115212
rect 265158 115200 265164 115212
rect 265216 115200 265222 115252
rect 166994 113772 167000 113824
rect 167052 113812 167058 113824
rect 265066 113812 265072 113824
rect 167052 113784 265072 113812
rect 167052 113772 167058 113784
rect 265066 113772 265072 113784
rect 265124 113772 265130 113824
rect 442258 113092 442264 113144
rect 442316 113132 442322 113144
rect 579798 113132 579804 113144
rect 442316 113104 579804 113132
rect 442316 113092 442322 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 173894 112412 173900 112464
rect 173952 112452 173958 112464
rect 266630 112452 266636 112464
rect 173952 112424 266636 112452
rect 173952 112412 173958 112424
rect 266630 112412 266636 112424
rect 266688 112412 266694 112464
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 86218 111772 86224 111784
rect 3200 111744 86224 111772
rect 3200 111732 3206 111744
rect 86218 111732 86224 111744
rect 86276 111732 86282 111784
rect 185026 111052 185032 111104
rect 185084 111092 185090 111104
rect 267734 111092 267740 111104
rect 185084 111064 267740 111092
rect 185084 111052 185090 111064
rect 267734 111052 267740 111064
rect 267792 111052 267798 111104
rect 269850 111052 269856 111104
rect 269908 111092 269914 111104
rect 280522 111092 280528 111104
rect 269908 111064 280528 111092
rect 269908 111052 269914 111064
rect 280522 111052 280528 111064
rect 280580 111052 280586 111104
rect 191834 109692 191840 109744
rect 191892 109732 191898 109744
rect 269298 109732 269304 109744
rect 191892 109704 269304 109732
rect 191892 109692 191898 109704
rect 269298 109692 269304 109704
rect 269356 109692 269362 109744
rect 131114 108264 131120 108316
rect 131172 108304 131178 108316
rect 259454 108304 259460 108316
rect 131172 108276 259460 108304
rect 131172 108264 131178 108276
rect 259454 108264 259460 108276
rect 259512 108264 259518 108316
rect 260098 108264 260104 108316
rect 260156 108304 260162 108316
rect 278958 108304 278964 108316
rect 260156 108276 278964 108304
rect 260156 108264 260162 108276
rect 278958 108264 278964 108276
rect 279016 108264 279022 108316
rect 201586 106904 201592 106956
rect 201644 106944 201650 106956
rect 270494 106944 270500 106956
rect 201644 106916 270500 106944
rect 201644 106904 201650 106916
rect 270494 106904 270500 106916
rect 270552 106904 270558 106956
rect 219434 105612 219440 105664
rect 219492 105652 219498 105664
rect 273254 105652 273260 105664
rect 219492 105624 273260 105652
rect 219492 105612 219498 105624
rect 273254 105612 273260 105624
rect 273312 105612 273318 105664
rect 124214 105544 124220 105596
rect 124272 105584 124278 105596
rect 258166 105584 258172 105596
rect 124272 105556 258172 105584
rect 124272 105544 124278 105556
rect 258166 105544 258172 105556
rect 258224 105544 258230 105596
rect 230474 104184 230480 104236
rect 230532 104224 230538 104236
rect 274726 104224 274732 104236
rect 230532 104196 274732 104224
rect 230532 104184 230538 104196
rect 274726 104184 274732 104196
rect 274784 104184 274790 104236
rect 106274 104116 106280 104168
rect 106332 104156 106338 104168
rect 255590 104156 255596 104168
rect 106332 104128 255596 104156
rect 106332 104116 106338 104128
rect 255590 104116 255596 104128
rect 255648 104116 255654 104168
rect 135346 102756 135352 102808
rect 135404 102796 135410 102808
rect 261018 102796 261024 102808
rect 135404 102768 261024 102796
rect 135404 102756 135410 102768
rect 261018 102756 261024 102768
rect 261076 102756 261082 102808
rect 138014 101396 138020 101448
rect 138072 101436 138078 101448
rect 260926 101436 260932 101448
rect 138072 101408 260932 101436
rect 138072 101396 138078 101408
rect 260926 101396 260932 101408
rect 260984 101396 260990 101448
rect 149054 99968 149060 100020
rect 149112 100008 149118 100020
rect 262766 100008 262772 100020
rect 149112 99980 262772 100008
rect 149112 99968 149118 99980
rect 262766 99968 262772 99980
rect 262824 99968 262830 100020
rect 151906 98608 151912 98660
rect 151964 98648 151970 98660
rect 263686 98648 263692 98660
rect 151964 98620 263692 98648
rect 151964 98608 151970 98620
rect 263686 98608 263692 98620
rect 263744 98608 263750 98660
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 10318 97968 10324 97980
rect 3568 97940 10324 97968
rect 3568 97928 3574 97940
rect 10318 97928 10324 97940
rect 10376 97928 10382 97980
rect 114554 95888 114560 95940
rect 114612 95928 114618 95940
rect 256878 95928 256884 95940
rect 114612 95900 256884 95928
rect 114612 95888 114618 95900
rect 256878 95888 256884 95900
rect 256936 95888 256942 95940
rect 4798 94460 4804 94512
rect 4856 94500 4862 94512
rect 238754 94500 238760 94512
rect 4856 94472 238760 94500
rect 4856 94460 4862 94472
rect 238754 94460 238760 94472
rect 238812 94460 238818 94512
rect 102134 93100 102140 93152
rect 102192 93140 102198 93152
rect 255498 93140 255504 93152
rect 102192 93112 255504 93140
rect 102192 93100 102198 93112
rect 255498 93100 255504 93112
rect 255556 93100 255562 93152
rect 111794 91740 111800 91792
rect 111852 91780 111858 91792
rect 256786 91780 256792 91792
rect 111852 91752 256792 91780
rect 111852 91740 111858 91752
rect 256786 91740 256792 91752
rect 256844 91740 256850 91792
rect 122834 90312 122840 90364
rect 122892 90352 122898 90364
rect 258534 90352 258540 90364
rect 122892 90324 258540 90352
rect 122892 90312 122898 90324
rect 258534 90312 258540 90324
rect 258592 90312 258598 90364
rect 241606 89224 241612 89276
rect 241664 89264 241670 89276
rect 277854 89264 277860 89276
rect 241664 89236 277860 89264
rect 241664 89224 241670 89236
rect 277854 89224 277860 89236
rect 277912 89224 277918 89276
rect 238754 89156 238760 89208
rect 238812 89196 238818 89208
rect 276198 89196 276204 89208
rect 238812 89168 276204 89196
rect 238812 89156 238818 89168
rect 276198 89156 276204 89168
rect 276256 89156 276262 89208
rect 235994 89088 236000 89140
rect 236052 89128 236058 89140
rect 276290 89128 276296 89140
rect 236052 89100 276296 89128
rect 236052 89088 236058 89100
rect 276290 89088 276296 89100
rect 276348 89088 276354 89140
rect 233234 89020 233240 89072
rect 233292 89060 233298 89072
rect 276382 89060 276388 89072
rect 233292 89032 276388 89060
rect 233292 89020 233298 89032
rect 276382 89020 276388 89032
rect 276440 89020 276446 89072
rect 290274 89020 290280 89072
rect 290332 89060 290338 89072
rect 322934 89060 322940 89072
rect 290332 89032 322940 89060
rect 290332 89020 290338 89032
rect 322934 89020 322940 89032
rect 322992 89020 322998 89072
rect 99374 88952 99380 89004
rect 99432 88992 99438 89004
rect 247770 88992 247776 89004
rect 99432 88964 247776 88992
rect 99432 88952 99438 88964
rect 247770 88952 247776 88964
rect 247828 88952 247834 89004
rect 255498 88952 255504 89004
rect 255556 88992 255562 89004
rect 278038 88992 278044 89004
rect 255556 88964 278044 88992
rect 255556 88952 255562 88964
rect 278038 88952 278044 88964
rect 278096 88952 278102 89004
rect 290182 88952 290188 89004
rect 290240 88992 290246 89004
rect 325694 88992 325700 89004
rect 290240 88964 325700 88992
rect 290240 88952 290246 88964
rect 325694 88952 325700 88964
rect 325752 88952 325758 89004
rect 278958 88748 278964 88800
rect 279016 88788 279022 88800
rect 283282 88788 283288 88800
rect 279016 88760 283288 88788
rect 279016 88748 279022 88760
rect 283282 88748 283288 88760
rect 283340 88748 283346 88800
rect 45554 87592 45560 87644
rect 45612 87632 45618 87644
rect 246390 87632 246396 87644
rect 45612 87604 246396 87632
rect 45612 87592 45618 87604
rect 246390 87592 246396 87604
rect 246448 87592 246454 87644
rect 117314 86232 117320 86284
rect 117372 86272 117378 86284
rect 238018 86272 238024 86284
rect 117372 86244 238024 86272
rect 117372 86232 117378 86244
rect 238018 86232 238024 86244
rect 238076 86232 238082 86284
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 95878 85524 95884 85536
rect 3568 85496 95884 85524
rect 3568 85484 3574 85496
rect 95878 85484 95884 85496
rect 95936 85484 95942 85536
rect 287054 51688 287060 51740
rect 287112 51728 287118 51740
rect 307846 51728 307852 51740
rect 287112 51700 307852 51728
rect 287112 51688 287118 51700
rect 307846 51688 307852 51700
rect 307904 51688 307910 51740
rect 494698 33056 494704 33108
rect 494756 33096 494762 33108
rect 580166 33096 580172 33108
rect 494756 33068 580172 33096
rect 494756 33056 494762 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 24854 28228 24860 28280
rect 24912 28268 24918 28280
rect 243262 28268 243268 28280
rect 24912 28240 243268 28268
rect 24912 28228 24918 28240
rect 243262 28228 243268 28240
rect 243320 28228 243326 28280
rect 113174 26868 113180 26920
rect 113232 26908 113238 26920
rect 257154 26908 257160 26920
rect 113232 26880 257160 26908
rect 113232 26868 113238 26880
rect 257154 26868 257160 26880
rect 257212 26868 257218 26920
rect 110506 25508 110512 25560
rect 110564 25548 110570 25560
rect 242158 25548 242164 25560
rect 110564 25520 242164 25548
rect 110564 25508 110570 25520
rect 242158 25508 242164 25520
rect 242216 25508 242222 25560
rect 102226 24080 102232 24132
rect 102284 24120 102290 24132
rect 247678 24120 247684 24132
rect 102284 24092 247684 24120
rect 102284 24080 102290 24092
rect 247678 24080 247684 24092
rect 247736 24080 247742 24132
rect 88334 22720 88340 22772
rect 88392 22760 88398 22772
rect 246298 22760 246304 22772
rect 88392 22732 246304 22760
rect 88392 22720 88398 22732
rect 246298 22720 246304 22732
rect 246356 22720 246362 22772
rect 247402 22720 247408 22772
rect 247460 22760 247466 22772
rect 277762 22760 277768 22772
rect 247460 22732 277768 22760
rect 247460 22720 247466 22732
rect 277762 22720 277768 22732
rect 277820 22720 277826 22772
rect 290090 22720 290096 22772
rect 290148 22760 290154 22772
rect 324314 22760 324320 22772
rect 290148 22732 324320 22760
rect 290148 22720 290154 22732
rect 324314 22720 324320 22732
rect 324372 22720 324378 22772
rect 160094 21360 160100 21412
rect 160152 21400 160158 21412
rect 264514 21400 264520 21412
rect 160152 21372 264520 21400
rect 160152 21360 160158 21372
rect 264514 21360 264520 21372
rect 264572 21360 264578 21412
rect 142154 19932 142160 19984
rect 142212 19972 142218 19984
rect 260834 19972 260840 19984
rect 142212 19944 260840 19972
rect 142212 19932 142218 19944
rect 260834 19932 260840 19944
rect 260892 19932 260898 19984
rect 212534 18572 212540 18624
rect 212592 18612 212598 18624
rect 271966 18612 271972 18624
rect 212592 18584 271972 18612
rect 212592 18572 212598 18584
rect 271966 18572 271972 18584
rect 272024 18572 272030 18624
rect 291194 18572 291200 18624
rect 291252 18612 291258 18624
rect 329834 18612 329840 18624
rect 291252 18584 329840 18612
rect 291252 18572 291258 18584
rect 329834 18572 329840 18584
rect 329892 18572 329898 18624
rect 267734 17280 267740 17332
rect 267792 17320 267798 17332
rect 281626 17320 281632 17332
rect 267792 17292 281632 17320
rect 267792 17280 267798 17292
rect 281626 17280 281632 17292
rect 281684 17280 281690 17332
rect 194594 17212 194600 17264
rect 194652 17252 194658 17264
rect 269206 17252 269212 17264
rect 194652 17224 269212 17252
rect 194652 17212 194658 17224
rect 269206 17212 269212 17224
rect 269264 17212 269270 17264
rect 259454 15852 259460 15904
rect 259512 15892 259518 15904
rect 279510 15892 279516 15904
rect 259512 15864 279516 15892
rect 259512 15852 259518 15864
rect 279510 15852 279516 15864
rect 279568 15852 279574 15904
rect 119890 14424 119896 14476
rect 119948 14464 119954 14476
rect 253198 14464 253204 14476
rect 119948 14436 253204 14464
rect 119948 14424 119954 14436
rect 253198 14424 253204 14436
rect 253256 14424 253262 14476
rect 256694 14424 256700 14476
rect 256752 14464 256758 14476
rect 278866 14464 278872 14476
rect 256752 14436 278872 14464
rect 256752 14424 256758 14436
rect 278866 14424 278872 14436
rect 278924 14424 278930 14476
rect 288526 14424 288532 14476
rect 288584 14464 288590 14476
rect 312170 14464 312176 14476
rect 288584 14436 312176 14464
rect 288584 14424 288590 14436
rect 312170 14424 312176 14436
rect 312228 14424 312234 14476
rect 109034 13064 109040 13116
rect 109092 13104 109098 13116
rect 255958 13104 255964 13116
rect 109092 13076 255964 13104
rect 109092 13064 109098 13076
rect 255958 13064 255964 13076
rect 256016 13064 256022 13116
rect 184934 11772 184940 11824
rect 184992 11812 184998 11824
rect 186130 11812 186136 11824
rect 184992 11784 186136 11812
rect 184992 11772 184998 11784
rect 186130 11772 186136 11784
rect 186188 11772 186194 11824
rect 105722 11704 105728 11756
rect 105780 11744 105786 11756
rect 255406 11744 255412 11756
rect 105780 11716 255412 11744
rect 105780 11704 105786 11716
rect 255406 11704 255412 11716
rect 255464 11704 255470 11756
rect 278038 11568 278044 11620
rect 278096 11608 278102 11620
rect 283190 11608 283196 11620
rect 278096 11580 283196 11608
rect 278096 11568 278102 11580
rect 283190 11568 283196 11580
rect 283248 11568 283254 11620
rect 227530 10344 227536 10396
rect 227588 10384 227594 10396
rect 275094 10384 275100 10396
rect 227588 10356 275100 10384
rect 227588 10344 227594 10356
rect 275094 10344 275100 10356
rect 275152 10344 275158 10396
rect 274818 10276 274824 10328
rect 274876 10316 274882 10328
rect 280798 10316 280804 10328
rect 274876 10288 280804 10316
rect 274876 10276 274882 10288
rect 280798 10276 280804 10288
rect 280856 10276 280862 10328
rect 298094 10276 298100 10328
rect 298152 10316 298158 10328
rect 376018 10316 376024 10328
rect 298152 10288 376024 10316
rect 298152 10276 298158 10288
rect 376018 10276 376024 10288
rect 376076 10276 376082 10328
rect 294598 9188 294604 9240
rect 294656 9228 294662 9240
rect 344554 9228 344560 9240
rect 294656 9200 344560 9228
rect 294656 9188 294662 9200
rect 344554 9188 344560 9200
rect 344612 9188 344618 9240
rect 294230 9120 294236 9172
rect 294288 9160 294294 9172
rect 348050 9160 348056 9172
rect 294288 9132 348056 9160
rect 294288 9120 294294 9132
rect 348050 9120 348056 9132
rect 348108 9120 348114 9172
rect 296070 9052 296076 9104
rect 296128 9092 296134 9104
rect 355226 9092 355232 9104
rect 296128 9064 355232 9092
rect 296128 9052 296134 9064
rect 355226 9052 355232 9064
rect 355284 9052 355290 9104
rect 299382 8984 299388 9036
rect 299440 9024 299446 9036
rect 397730 9024 397736 9036
rect 299440 8996 397736 9024
rect 299440 8984 299446 8996
rect 397730 8984 397736 8996
rect 397788 8984 397794 9036
rect 87966 8916 87972 8968
rect 88024 8956 88030 8968
rect 252922 8956 252928 8968
rect 88024 8928 252928 8956
rect 88024 8916 88030 8928
rect 252922 8916 252928 8928
rect 252980 8916 252986 8968
rect 284662 8916 284668 8968
rect 284720 8956 284726 8968
rect 292482 8956 292488 8968
rect 284720 8928 292488 8956
rect 284720 8916 284726 8928
rect 292482 8916 292488 8928
rect 292540 8916 292546 8968
rect 295058 8916 295064 8968
rect 295116 8956 295122 8968
rect 414290 8956 414296 8968
rect 295116 8928 414296 8956
rect 295116 8916 295122 8928
rect 414290 8916 414296 8928
rect 414348 8916 414354 8968
rect 177850 7624 177856 7676
rect 177908 7664 177914 7676
rect 266538 7664 266544 7676
rect 177908 7636 266544 7664
rect 177908 7624 177914 7636
rect 266538 7624 266544 7636
rect 266596 7624 266602 7676
rect 295518 7624 295524 7676
rect 295576 7664 295582 7676
rect 295576 7636 302234 7664
rect 295576 7624 295582 7636
rect 39574 7556 39580 7608
rect 39632 7596 39638 7608
rect 246022 7596 246028 7608
rect 39632 7568 246028 7596
rect 39632 7556 39638 7568
rect 246022 7556 246028 7568
rect 246080 7556 246086 7608
rect 299566 7556 299572 7608
rect 299624 7596 299630 7608
rect 300762 7596 300768 7608
rect 299624 7568 300768 7596
rect 299624 7556 299630 7568
rect 300762 7556 300768 7568
rect 300820 7556 300826 7608
rect 302206 7596 302234 7636
rect 361114 7596 361120 7608
rect 302206 7568 361120 7596
rect 361114 7556 361120 7568
rect 361172 7556 361178 7608
rect 261754 6876 261760 6928
rect 261812 6916 261818 6928
rect 269758 6916 269764 6928
rect 261812 6888 269764 6916
rect 261812 6876 261818 6888
rect 269758 6876 269764 6888
rect 269816 6876 269822 6928
rect 284570 6876 284576 6928
rect 284628 6916 284634 6928
rect 288986 6916 288992 6928
rect 284628 6888 288992 6916
rect 284628 6876 284634 6888
rect 288986 6876 288992 6888
rect 289044 6876 289050 6928
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 14458 6848 14464 6860
rect 3476 6820 14464 6848
rect 3476 6808 3482 6820
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 288434 6808 288440 6860
rect 288492 6848 288498 6860
rect 316218 6848 316224 6860
rect 288492 6820 316224 6848
rect 288492 6808 288498 6820
rect 316218 6808 316224 6820
rect 316276 6808 316282 6860
rect 289998 6740 290004 6792
rect 290056 6780 290062 6792
rect 322106 6780 322112 6792
rect 290056 6752 322112 6780
rect 290056 6740 290062 6752
rect 322106 6740 322112 6752
rect 322164 6740 322170 6792
rect 242894 6672 242900 6724
rect 242952 6712 242958 6724
rect 277670 6712 277676 6724
rect 242952 6684 277676 6712
rect 242952 6672 242958 6684
rect 277670 6672 277676 6684
rect 277728 6672 277734 6724
rect 294138 6672 294144 6724
rect 294196 6712 294202 6724
rect 350442 6712 350448 6724
rect 294196 6684 350448 6712
rect 294196 6672 294202 6684
rect 350442 6672 350448 6684
rect 350500 6672 350506 6724
rect 234614 6604 234620 6656
rect 234672 6644 234678 6656
rect 276566 6644 276572 6656
rect 234672 6616 276572 6644
rect 234672 6604 234678 6616
rect 276566 6604 276572 6616
rect 276624 6604 276630 6656
rect 294046 6604 294052 6656
rect 294104 6644 294110 6656
rect 354030 6644 354036 6656
rect 294104 6616 354036 6644
rect 294104 6604 294110 6616
rect 354030 6604 354036 6616
rect 354088 6604 354094 6656
rect 235810 6536 235816 6588
rect 235868 6576 235874 6588
rect 276106 6576 276112 6588
rect 235868 6548 276112 6576
rect 235868 6536 235874 6548
rect 276106 6536 276112 6548
rect 276164 6536 276170 6588
rect 295426 6536 295432 6588
rect 295484 6576 295490 6588
rect 357526 6576 357532 6588
rect 295484 6548 357532 6576
rect 295484 6536 295490 6548
rect 357526 6536 357532 6548
rect 357584 6536 357590 6588
rect 176654 6468 176660 6520
rect 176712 6508 176718 6520
rect 257338 6508 257344 6520
rect 176712 6480 257344 6508
rect 176712 6468 176718 6480
rect 257338 6468 257344 6480
rect 257396 6468 257402 6520
rect 285766 6468 285772 6520
rect 285824 6508 285830 6520
rect 294874 6508 294880 6520
rect 285824 6480 294880 6508
rect 285824 6468 285830 6480
rect 294874 6468 294880 6480
rect 294932 6468 294938 6520
rect 296714 6468 296720 6520
rect 296772 6508 296778 6520
rect 365806 6508 365812 6520
rect 296772 6480 365812 6508
rect 296772 6468 296778 6480
rect 365806 6468 365812 6480
rect 365864 6468 365870 6520
rect 173158 6400 173164 6452
rect 173216 6440 173222 6452
rect 266446 6440 266452 6452
rect 173216 6412 266452 6440
rect 173216 6400 173222 6412
rect 266446 6400 266452 6412
rect 266504 6400 266510 6452
rect 290642 6400 290648 6452
rect 290700 6440 290706 6452
rect 400122 6440 400128 6452
rect 290700 6412 400128 6440
rect 290700 6400 290706 6412
rect 400122 6400 400128 6412
rect 400180 6400 400186 6452
rect 101030 6332 101036 6384
rect 101088 6372 101094 6384
rect 255774 6372 255780 6384
rect 101088 6344 255780 6372
rect 101088 6332 101094 6344
rect 255774 6332 255780 6344
rect 255832 6332 255838 6384
rect 286962 6332 286968 6384
rect 287020 6372 287026 6384
rect 403618 6372 403624 6384
rect 287020 6344 403624 6372
rect 287020 6332 287026 6344
rect 403618 6332 403624 6344
rect 403676 6332 403682 6384
rect 70302 6264 70308 6316
rect 70360 6304 70366 6316
rect 250254 6304 250260 6316
rect 70360 6276 250260 6304
rect 70360 6264 70366 6276
rect 250254 6264 250260 6276
rect 250312 6264 250318 6316
rect 293586 6264 293592 6316
rect 293644 6304 293650 6316
rect 410794 6304 410800 6316
rect 293644 6276 410800 6304
rect 293644 6264 293650 6276
rect 410794 6264 410800 6276
rect 410852 6264 410858 6316
rect 52546 6196 52552 6248
rect 52604 6236 52610 6248
rect 247310 6236 247316 6248
rect 52604 6208 247316 6236
rect 52604 6196 52610 6208
rect 247310 6196 247316 6208
rect 247368 6196 247374 6248
rect 254670 6196 254676 6248
rect 254728 6236 254734 6248
rect 279234 6236 279240 6248
rect 254728 6208 279240 6236
rect 254728 6196 254734 6208
rect 279234 6196 279240 6208
rect 279292 6196 279298 6248
rect 289722 6196 289728 6248
rect 289780 6236 289786 6248
rect 408402 6236 408408 6248
rect 289780 6208 408408 6236
rect 289780 6196 289786 6208
rect 408402 6196 408408 6208
rect 408460 6196 408466 6248
rect 45462 6128 45468 6180
rect 45520 6168 45526 6180
rect 244918 6168 244924 6180
rect 45520 6140 244924 6168
rect 45520 6128 45526 6140
rect 244918 6128 244924 6140
rect 244976 6128 244982 6180
rect 248782 6128 248788 6180
rect 248840 6168 248846 6180
rect 277578 6168 277584 6180
rect 248840 6140 277584 6168
rect 248840 6128 248846 6140
rect 277578 6128 277584 6140
rect 277636 6128 277642 6180
rect 288342 6128 288348 6180
rect 288400 6168 288406 6180
rect 407206 6168 407212 6180
rect 288400 6140 407212 6168
rect 288400 6128 288406 6140
rect 407206 6128 407212 6140
rect 407264 6128 407270 6180
rect 293310 5448 293316 5500
rect 293368 5488 293374 5500
rect 297266 5488 297272 5500
rect 293368 5460 297272 5488
rect 293368 5448 293374 5460
rect 297266 5448 297272 5460
rect 297324 5448 297330 5500
rect 210970 5244 210976 5296
rect 211028 5284 211034 5296
rect 268378 5284 268384 5296
rect 211028 5256 268384 5284
rect 211028 5244 211034 5256
rect 268378 5244 268384 5256
rect 268436 5244 268442 5296
rect 207382 5176 207388 5228
rect 207440 5216 207446 5228
rect 272426 5216 272432 5228
rect 207440 5188 272432 5216
rect 207440 5176 207446 5188
rect 272426 5176 272432 5188
rect 272484 5176 272490 5228
rect 297358 5176 297364 5228
rect 297416 5216 297422 5228
rect 297416 5188 302234 5216
rect 297416 5176 297422 5188
rect 189718 5108 189724 5160
rect 189776 5148 189782 5160
rect 269942 5148 269948 5160
rect 189776 5120 269948 5148
rect 189776 5108 189782 5120
rect 269942 5108 269948 5120
rect 270000 5108 270006 5160
rect 289814 5108 289820 5160
rect 289872 5148 289878 5160
rect 289872 5120 298692 5148
rect 289872 5108 289878 5120
rect 169570 5040 169576 5092
rect 169628 5080 169634 5092
rect 266906 5080 266912 5092
rect 169628 5052 266912 5080
rect 169628 5040 169634 5052
rect 266906 5040 266912 5052
rect 266964 5040 266970 5092
rect 285674 5040 285680 5092
rect 285732 5080 285738 5092
rect 298462 5080 298468 5092
rect 285732 5052 298468 5080
rect 285732 5040 285738 5052
rect 298462 5040 298468 5052
rect 298520 5040 298526 5092
rect 164878 4972 164884 5024
rect 164936 5012 164942 5024
rect 265526 5012 265532 5024
rect 164936 4984 265532 5012
rect 164936 4972 164942 4984
rect 265526 4972 265532 4984
rect 265584 4972 265590 5024
rect 289906 4972 289912 5024
rect 289964 5012 289970 5024
rect 297358 5012 297364 5024
rect 289964 4984 297364 5012
rect 289964 4972 289970 4984
rect 297358 4972 297364 4984
rect 297416 4972 297422 5024
rect 97442 4904 97448 4956
rect 97500 4944 97506 4956
rect 254118 4944 254124 4956
rect 97500 4916 254124 4944
rect 97500 4904 97506 4916
rect 254118 4904 254124 4916
rect 254176 4904 254182 4956
rect 265342 4904 265348 4956
rect 265400 4944 265406 4956
rect 279418 4944 279424 4956
rect 265400 4916 279424 4944
rect 265400 4904 265406 4916
rect 279418 4904 279424 4916
rect 279476 4904 279482 4956
rect 298664 4944 298692 5120
rect 302206 5080 302234 5188
rect 327994 5080 328000 5092
rect 302206 5052 306374 5080
rect 306346 5012 306374 5052
rect 325666 5052 328000 5080
rect 324406 5012 324412 5024
rect 306346 4984 324412 5012
rect 324406 4972 324412 4984
rect 324464 4972 324470 5024
rect 325666 4944 325694 5052
rect 327994 5040 328000 5052
rect 328052 5040 328058 5092
rect 298664 4916 325694 4944
rect 48958 4836 48964 4888
rect 49016 4876 49022 4888
rect 247218 4876 247224 4888
rect 49016 4848 247224 4876
rect 49016 4836 49022 4848
rect 247218 4836 247224 4848
rect 247276 4836 247282 4888
rect 277486 4876 277492 4888
rect 272536 4848 277492 4876
rect 15930 4768 15936 4820
rect 15988 4808 15994 4820
rect 241974 4808 241980 4820
rect 15988 4780 241980 4808
rect 15988 4768 15994 4780
rect 241974 4768 241980 4780
rect 242032 4768 242038 4820
rect 245194 4768 245200 4820
rect 245252 4808 245258 4820
rect 272536 4808 272564 4848
rect 277486 4836 277492 4848
rect 277544 4836 277550 4888
rect 293954 4836 293960 4888
rect 294012 4876 294018 4888
rect 349246 4876 349252 4888
rect 294012 4848 349252 4876
rect 294012 4836 294018 4848
rect 349246 4836 349252 4848
rect 349304 4836 349310 4888
rect 245252 4780 272564 4808
rect 245252 4768 245258 4780
rect 295334 4768 295340 4820
rect 295392 4808 295398 4820
rect 359918 4808 359924 4820
rect 295392 4780 359924 4808
rect 295392 4768 295398 4780
rect 359918 4768 359924 4780
rect 359976 4768 359982 4820
rect 278682 4360 278688 4412
rect 278740 4400 278746 4412
rect 282086 4400 282092 4412
rect 278740 4372 282092 4400
rect 278740 4360 278746 4372
rect 282086 4360 282092 4372
rect 282144 4360 282150 4412
rect 287698 4156 287704 4208
rect 287756 4196 287762 4208
rect 290182 4196 290188 4208
rect 287756 4168 290188 4196
rect 287756 4156 287762 4168
rect 290182 4156 290188 4168
rect 290240 4156 290246 4208
rect 12342 4088 12348 4140
rect 12400 4128 12406 4140
rect 18598 4128 18604 4140
rect 12400 4100 18604 4128
rect 12400 4088 12406 4100
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 253474 4088 253480 4140
rect 253532 4128 253538 4140
rect 260190 4128 260196 4140
rect 253532 4100 260196 4128
rect 253532 4088 253538 4100
rect 260190 4088 260196 4100
rect 260248 4088 260254 4140
rect 285582 4088 285588 4140
rect 285640 4128 285646 4140
rect 338666 4128 338672 4140
rect 285640 4100 338672 4128
rect 285640 4088 285646 4100
rect 338666 4088 338672 4100
rect 338724 4088 338730 4140
rect 429654 4088 429660 4140
rect 429712 4128 429718 4140
rect 440510 4128 440516 4140
rect 429712 4100 440516 4128
rect 429712 4088 429718 4100
rect 440510 4088 440516 4100
rect 440568 4088 440574 4140
rect 292390 4020 292396 4072
rect 292448 4060 292454 4072
rect 297450 4060 297456 4072
rect 292448 4032 297456 4060
rect 292448 4020 292454 4032
rect 297450 4020 297456 4032
rect 297508 4020 297514 4072
rect 298738 4020 298744 4072
rect 298796 4060 298802 4072
rect 369394 4060 369400 4072
rect 298796 4032 369400 4060
rect 298796 4020 298802 4032
rect 369394 4020 369400 4032
rect 369452 4020 369458 4072
rect 427262 4020 427268 4072
rect 427320 4060 427326 4072
rect 437842 4060 437848 4072
rect 427320 4032 437848 4060
rect 427320 4020 427326 4032
rect 437842 4020 437848 4032
rect 437900 4020 437906 4072
rect 6454 3952 6460 4004
rect 6512 3992 6518 4004
rect 7650 3992 7656 4004
rect 6512 3964 7656 3992
rect 6512 3952 6518 3964
rect 7650 3952 7656 3964
rect 7708 3952 7714 4004
rect 295242 3952 295248 4004
rect 295300 3992 295306 4004
rect 384758 3992 384764 4004
rect 295300 3964 384764 3992
rect 295300 3952 295306 3964
rect 384758 3952 384764 3964
rect 384816 3952 384822 4004
rect 426158 3952 426164 4004
rect 426216 3992 426222 4004
rect 437474 3992 437480 4004
rect 426216 3964 437480 3992
rect 426216 3952 426222 3964
rect 437474 3952 437480 3964
rect 437532 3952 437538 4004
rect 266538 3884 266544 3936
rect 266596 3924 266602 3936
rect 269850 3924 269856 3936
rect 266596 3896 269856 3924
rect 266596 3884 266602 3896
rect 269850 3884 269856 3896
rect 269908 3884 269914 3936
rect 293862 3884 293868 3936
rect 293920 3924 293926 3936
rect 391842 3924 391848 3936
rect 293920 3896 391848 3924
rect 293920 3884 293926 3896
rect 391842 3884 391848 3896
rect 391900 3884 391906 3936
rect 423766 3884 423772 3936
rect 423824 3924 423830 3936
rect 437658 3924 437664 3936
rect 423824 3896 437664 3924
rect 423824 3884 423830 3896
rect 437658 3884 437664 3896
rect 437716 3884 437722 3936
rect 5258 3816 5264 3868
rect 5316 3856 5322 3868
rect 7558 3856 7564 3868
rect 5316 3828 7564 3856
rect 5316 3816 5322 3828
rect 7558 3816 7564 3828
rect 7616 3816 7622 3868
rect 171962 3816 171968 3868
rect 172020 3856 172026 3868
rect 239398 3856 239404 3868
rect 172020 3828 239404 3856
rect 172020 3816 172026 3828
rect 239398 3816 239404 3828
rect 239456 3816 239462 3868
rect 293770 3816 293776 3868
rect 293828 3856 293834 3868
rect 395338 3856 395344 3868
rect 293828 3828 395344 3856
rect 293828 3816 293834 3828
rect 395338 3816 395344 3828
rect 395396 3816 395402 3868
rect 424962 3816 424968 3868
rect 425020 3856 425026 3868
rect 439130 3856 439136 3868
rect 425020 3828 439136 3856
rect 425020 3816 425026 3828
rect 439130 3816 439136 3828
rect 439188 3816 439194 3868
rect 460198 3816 460204 3868
rect 460256 3856 460262 3868
rect 462774 3856 462780 3868
rect 460256 3828 462780 3856
rect 460256 3816 460262 3828
rect 462774 3816 462780 3828
rect 462832 3816 462838 3868
rect 516778 3816 516784 3868
rect 516836 3856 516842 3868
rect 519538 3856 519544 3868
rect 516836 3828 519544 3856
rect 516836 3816 516842 3828
rect 519538 3816 519544 3828
rect 519596 3816 519602 3868
rect 566458 3816 566464 3868
rect 566516 3856 566522 3868
rect 569126 3856 569132 3868
rect 566516 3828 569132 3856
rect 566516 3816 566522 3828
rect 569126 3816 569132 3828
rect 569184 3816 569190 3868
rect 135254 3748 135260 3800
rect 135312 3788 135318 3800
rect 136450 3788 136456 3800
rect 135312 3760 136456 3788
rect 135312 3748 135318 3760
rect 136450 3748 136456 3760
rect 136508 3748 136514 3800
rect 161290 3748 161296 3800
rect 161348 3788 161354 3800
rect 264238 3788 264244 3800
rect 161348 3760 264244 3788
rect 161348 3748 161354 3760
rect 264238 3748 264244 3760
rect 264296 3748 264302 3800
rect 294966 3748 294972 3800
rect 295024 3788 295030 3800
rect 295024 3760 298048 3788
rect 295024 3748 295030 3760
rect 125870 3680 125876 3732
rect 125928 3720 125934 3732
rect 238110 3720 238116 3732
rect 125928 3692 238116 3720
rect 125928 3680 125934 3692
rect 238110 3680 238116 3692
rect 238168 3680 238174 3732
rect 244090 3680 244096 3732
rect 244148 3720 244154 3732
rect 278130 3720 278136 3732
rect 244148 3692 278136 3720
rect 244148 3680 244154 3692
rect 278130 3680 278136 3692
rect 278188 3680 278194 3732
rect 296622 3680 296628 3732
rect 296680 3720 296686 3732
rect 298020 3720 298048 3760
rect 298094 3748 298100 3800
rect 298152 3788 298158 3800
rect 398926 3788 398932 3800
rect 298152 3760 398932 3788
rect 298152 3748 298158 3760
rect 398926 3748 398932 3760
rect 398984 3748 398990 3800
rect 422570 3748 422576 3800
rect 422628 3788 422634 3800
rect 438946 3788 438952 3800
rect 422628 3760 438952 3788
rect 422628 3748 422634 3760
rect 438946 3748 438952 3760
rect 439004 3748 439010 3800
rect 402514 3720 402520 3732
rect 296680 3692 297588 3720
rect 298020 3692 402520 3720
rect 296680 3680 296686 3692
rect 13078 3652 13084 3664
rect 6886 3624 13084 3652
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 6886 3584 6914 3624
rect 13078 3612 13084 3624
rect 13136 3612 13142 3664
rect 28902 3612 28908 3664
rect 28960 3652 28966 3664
rect 39298 3652 39304 3664
rect 28960 3624 39304 3652
rect 28960 3612 28966 3624
rect 39298 3612 39304 3624
rect 39356 3612 39362 3664
rect 43070 3612 43076 3664
rect 43128 3652 43134 3664
rect 57238 3652 57244 3664
rect 43128 3624 57244 3652
rect 43128 3612 43134 3624
rect 57238 3612 57244 3624
rect 57296 3612 57302 3664
rect 68278 3652 68284 3664
rect 64846 3624 68284 3652
rect 2924 3556 6914 3584
rect 2924 3544 2930 3556
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 7708 3556 16574 3584
rect 7708 3544 7714 3556
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 4798 3516 4804 3528
rect 624 3488 4804 3516
rect 624 3476 630 3488
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 11698 3516 11704 3528
rect 10008 3488 11704 3516
rect 10008 3476 10014 3488
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 16546 3516 16574 3556
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 64846 3584 64874 3624
rect 68278 3612 68284 3624
rect 68336 3612 68342 3664
rect 93946 3612 93952 3664
rect 94004 3652 94010 3664
rect 254394 3652 254400 3664
rect 94004 3624 254400 3652
rect 94004 3612 94010 3624
rect 254394 3612 254400 3624
rect 254452 3612 254458 3664
rect 264146 3612 264152 3664
rect 264204 3652 264210 3664
rect 273898 3652 273904 3664
rect 264204 3624 273904 3652
rect 264204 3612 264210 3624
rect 273898 3612 273904 3624
rect 273956 3612 273962 3664
rect 291102 3612 291108 3664
rect 291160 3652 291166 3664
rect 297560 3652 297588 3692
rect 402514 3680 402520 3692
rect 402572 3680 402578 3732
rect 421374 3680 421380 3732
rect 421432 3720 421438 3732
rect 438026 3720 438032 3732
rect 421432 3692 438032 3720
rect 421432 3680 421438 3692
rect 438026 3680 438032 3692
rect 438084 3680 438090 3732
rect 409598 3652 409604 3664
rect 291160 3624 297404 3652
rect 297560 3624 409604 3652
rect 291160 3612 291166 3624
rect 20680 3556 64874 3584
rect 20680 3544 20686 3556
rect 67910 3544 67916 3596
rect 67968 3584 67974 3596
rect 71038 3584 71044 3596
rect 67968 3556 71044 3584
rect 67968 3544 67974 3556
rect 71038 3544 71044 3556
rect 71096 3544 71102 3596
rect 77294 3544 77300 3596
rect 77352 3584 77358 3596
rect 78214 3584 78220 3596
rect 77352 3556 78220 3584
rect 77352 3544 77358 3556
rect 78214 3544 78220 3556
rect 78272 3544 78278 3596
rect 85666 3544 85672 3596
rect 85724 3584 85730 3596
rect 88978 3584 88984 3596
rect 85724 3556 88984 3584
rect 85724 3544 85730 3556
rect 88978 3544 88984 3556
rect 89036 3544 89042 3596
rect 90358 3544 90364 3596
rect 90416 3584 90422 3596
rect 254302 3584 254308 3596
rect 90416 3556 254308 3584
rect 90416 3544 90422 3556
rect 254302 3544 254308 3556
rect 254360 3544 254366 3596
rect 262950 3544 262956 3596
rect 263008 3584 263014 3596
rect 266998 3584 267004 3596
rect 263008 3556 267004 3584
rect 263008 3544 263014 3556
rect 266998 3544 267004 3556
rect 267056 3544 267062 3596
rect 267090 3544 267096 3596
rect 267148 3584 267154 3596
rect 271230 3584 271236 3596
rect 267148 3556 271236 3584
rect 267148 3544 267154 3556
rect 271230 3544 271236 3556
rect 271288 3544 271294 3596
rect 283006 3544 283012 3596
rect 283064 3544 283070 3596
rect 284294 3544 284300 3596
rect 284352 3584 284358 3596
rect 285030 3584 285036 3596
rect 284352 3556 285036 3584
rect 284352 3544 284358 3556
rect 285030 3544 285036 3556
rect 285088 3544 285094 3596
rect 17218 3516 17224 3528
rect 16546 3488 17224 3516
rect 17218 3476 17224 3488
rect 17276 3476 17282 3528
rect 21818 3476 21824 3528
rect 21876 3516 21882 3528
rect 22738 3516 22744 3528
rect 21876 3488 22744 3516
rect 21876 3476 21882 3488
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24268 3488 29316 3516
rect 24268 3476 24274 3488
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 4890 3448 4896 3460
rect 4120 3420 4896 3448
rect 4120 3408 4126 3420
rect 4890 3408 4896 3420
rect 4948 3408 4954 3460
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 29288 3448 29316 3488
rect 30098 3476 30104 3528
rect 30156 3516 30162 3528
rect 31018 3516 31024 3528
rect 30156 3488 31024 3516
rect 30156 3476 30162 3488
rect 31018 3476 31024 3488
rect 31076 3476 31082 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 35158 3516 35164 3528
rect 33652 3488 35164 3516
rect 33652 3476 33658 3488
rect 35158 3476 35164 3488
rect 35216 3476 35222 3528
rect 38378 3476 38384 3528
rect 38436 3516 38442 3528
rect 39390 3516 39396 3528
rect 38436 3488 39396 3516
rect 38436 3476 38442 3488
rect 39390 3476 39396 3488
rect 39448 3476 39454 3528
rect 51350 3476 51356 3528
rect 51408 3516 51414 3528
rect 247678 3516 247684 3528
rect 51408 3488 247684 3516
rect 51408 3476 51414 3488
rect 247678 3476 247684 3488
rect 247736 3476 247742 3528
rect 251174 3476 251180 3528
rect 251232 3516 251238 3528
rect 268562 3516 268568 3528
rect 251232 3488 268568 3516
rect 251232 3476 251238 3488
rect 268562 3476 268568 3488
rect 268620 3476 268626 3528
rect 268838 3476 268844 3528
rect 268896 3516 268902 3528
rect 274082 3516 274088 3528
rect 268896 3488 274088 3516
rect 268896 3476 268902 3488
rect 274082 3476 274088 3488
rect 274140 3476 274146 3528
rect 277118 3476 277124 3528
rect 277176 3516 277182 3528
rect 282178 3516 282184 3528
rect 277176 3488 282184 3516
rect 277176 3476 277182 3488
rect 282178 3476 282184 3488
rect 282236 3476 282242 3528
rect 32398 3448 32404 3460
rect 11204 3420 26234 3448
rect 29288 3420 32404 3448
rect 11204 3408 11210 3420
rect 26206 3380 26234 3420
rect 32398 3408 32404 3420
rect 32456 3408 32462 3460
rect 35986 3408 35992 3460
rect 36044 3448 36050 3460
rect 50338 3448 50344 3460
rect 36044 3420 50344 3448
rect 36044 3408 36050 3420
rect 50338 3408 50344 3420
rect 50396 3408 50402 3460
rect 247126 3448 247132 3460
rect 55186 3420 247132 3448
rect 43438 3380 43444 3392
rect 26206 3352 43444 3380
rect 43438 3340 43444 3352
rect 43496 3340 43502 3392
rect 47854 3340 47860 3392
rect 47912 3380 47918 3392
rect 55186 3380 55214 3420
rect 247126 3408 247132 3420
rect 247184 3408 247190 3460
rect 249978 3408 249984 3460
rect 250036 3448 250042 3460
rect 268470 3448 268476 3460
rect 250036 3420 268476 3448
rect 250036 3408 250042 3420
rect 268470 3408 268476 3420
rect 268528 3408 268534 3460
rect 270034 3408 270040 3460
rect 270092 3448 270098 3460
rect 273990 3448 273996 3460
rect 270092 3420 273996 3448
rect 270092 3408 270098 3420
rect 273990 3408 273996 3420
rect 274048 3408 274054 3460
rect 276014 3408 276020 3460
rect 276072 3448 276078 3460
rect 283024 3448 283052 3544
rect 291838 3476 291844 3528
rect 291896 3516 291902 3528
rect 296070 3516 296076 3528
rect 291896 3488 296076 3516
rect 291896 3476 291902 3488
rect 296070 3476 296076 3488
rect 296128 3476 296134 3528
rect 297376 3516 297404 3624
rect 409598 3612 409604 3624
rect 409656 3612 409662 3664
rect 420178 3612 420184 3664
rect 420236 3652 420242 3664
rect 438854 3652 438860 3664
rect 420236 3624 438860 3652
rect 420236 3612 420242 3624
rect 438854 3612 438860 3624
rect 438912 3612 438918 3664
rect 297450 3544 297456 3596
rect 297508 3584 297514 3596
rect 406010 3584 406016 3596
rect 297508 3556 406016 3584
rect 297508 3544 297514 3556
rect 406010 3544 406016 3556
rect 406068 3544 406074 3596
rect 418982 3544 418988 3596
rect 419040 3584 419046 3596
rect 437566 3584 437572 3596
rect 419040 3556 437572 3584
rect 419040 3544 419046 3556
rect 437566 3544 437572 3556
rect 437624 3544 437630 3596
rect 442350 3544 442356 3596
rect 442408 3584 442414 3596
rect 447410 3584 447416 3596
rect 442408 3556 447416 3584
rect 442408 3544 442414 3556
rect 447410 3544 447416 3556
rect 447468 3544 447474 3596
rect 453298 3544 453304 3596
rect 453356 3584 453362 3596
rect 455690 3584 455696 3596
rect 453356 3556 455696 3584
rect 453356 3544 453362 3556
rect 455690 3544 455696 3556
rect 455748 3544 455754 3596
rect 467098 3544 467104 3596
rect 467156 3584 467162 3596
rect 469858 3584 469864 3596
rect 467156 3556 469864 3584
rect 467156 3544 467162 3556
rect 469858 3544 469864 3556
rect 469916 3544 469922 3596
rect 475378 3544 475384 3596
rect 475436 3584 475442 3596
rect 476942 3584 476948 3596
rect 475436 3556 476948 3584
rect 475436 3544 475442 3556
rect 476942 3544 476948 3556
rect 477000 3544 477006 3596
rect 500218 3544 500224 3596
rect 500276 3584 500282 3596
rect 501782 3584 501788 3596
rect 500276 3556 501788 3584
rect 500276 3544 500282 3556
rect 501782 3544 501788 3556
rect 501840 3544 501846 3596
rect 511258 3544 511264 3596
rect 511316 3584 511322 3596
rect 513558 3584 513564 3596
rect 511316 3556 513564 3584
rect 511316 3544 511322 3556
rect 513558 3544 513564 3556
rect 513616 3544 513622 3596
rect 413094 3516 413100 3528
rect 297376 3488 413100 3516
rect 413094 3476 413100 3488
rect 413152 3476 413158 3528
rect 417878 3476 417884 3528
rect 417936 3516 417942 3528
rect 439222 3516 439228 3528
rect 417936 3488 439228 3516
rect 417936 3476 417942 3488
rect 439222 3476 439228 3488
rect 439280 3476 439286 3528
rect 440326 3476 440332 3528
rect 440384 3516 440390 3528
rect 441522 3516 441528 3528
rect 440384 3488 441528 3516
rect 440384 3476 440390 3488
rect 441522 3476 441528 3488
rect 441580 3476 441586 3528
rect 448606 3476 448612 3528
rect 448664 3516 448670 3528
rect 449802 3516 449808 3528
rect 448664 3488 449808 3516
rect 448664 3476 448670 3488
rect 449802 3476 449808 3488
rect 449860 3476 449866 3528
rect 462958 3476 462964 3528
rect 463016 3516 463022 3528
rect 465166 3516 465172 3528
rect 463016 3488 465172 3516
rect 463016 3476 463022 3488
rect 465166 3476 465172 3488
rect 465224 3476 465230 3528
rect 538858 3476 538864 3528
rect 538916 3516 538922 3528
rect 540790 3516 540796 3528
rect 538916 3488 540796 3516
rect 538916 3476 538922 3488
rect 540790 3476 540796 3488
rect 540848 3476 540854 3528
rect 547874 3476 547880 3528
rect 547932 3516 547938 3528
rect 548702 3516 548708 3528
rect 547932 3488 548708 3516
rect 547932 3476 547938 3488
rect 548702 3476 548708 3488
rect 548760 3476 548766 3528
rect 556154 3476 556160 3528
rect 556212 3516 556218 3528
rect 556982 3516 556988 3528
rect 556212 3488 556988 3516
rect 556212 3476 556218 3488
rect 556982 3476 556988 3488
rect 557040 3476 557046 3528
rect 563698 3476 563704 3528
rect 563756 3516 563762 3528
rect 565630 3516 565636 3528
rect 563756 3488 565636 3516
rect 563756 3476 563762 3488
rect 565630 3476 565636 3488
rect 565688 3476 565694 3528
rect 571978 3476 571984 3528
rect 572036 3516 572042 3528
rect 573910 3516 573916 3528
rect 572036 3488 573916 3516
rect 572036 3476 572042 3488
rect 573910 3476 573916 3488
rect 573968 3476 573974 3528
rect 580994 3476 581000 3528
rect 581052 3516 581058 3528
rect 581822 3516 581828 3528
rect 581052 3488 581828 3516
rect 581052 3476 581058 3488
rect 581822 3476 581828 3488
rect 581880 3476 581886 3528
rect 276072 3420 283052 3448
rect 276072 3408 276078 3420
rect 292298 3408 292304 3460
rect 292356 3448 292362 3460
rect 416682 3448 416688 3460
rect 292356 3420 416688 3448
rect 292356 3408 292362 3420
rect 416682 3408 416688 3420
rect 416740 3408 416746 3460
rect 439038 3448 439044 3460
rect 422266 3420 439044 3448
rect 47912 3352 55214 3380
rect 47912 3340 47918 3352
rect 60734 3340 60740 3392
rect 60792 3380 60798 3392
rect 61654 3380 61660 3392
rect 60792 3352 61660 3380
rect 60792 3340 60798 3352
rect 61654 3340 61660 3352
rect 61712 3340 61718 3392
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 260650 3340 260656 3392
rect 260708 3380 260714 3392
rect 267090 3380 267096 3392
rect 260708 3352 267096 3380
rect 260708 3340 260714 3352
rect 267090 3340 267096 3352
rect 267148 3340 267154 3392
rect 295978 3340 295984 3392
rect 296036 3380 296042 3392
rect 346946 3380 346952 3392
rect 296036 3352 346952 3380
rect 296036 3340 296042 3352
rect 346946 3340 346952 3352
rect 347004 3340 347010 3392
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 358722 3380 358728 3392
rect 357492 3352 358728 3380
rect 357492 3340 357498 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 415486 3340 415492 3392
rect 415544 3380 415550 3392
rect 422266 3380 422294 3420
rect 439038 3408 439044 3420
rect 439096 3408 439102 3460
rect 445110 3408 445116 3460
rect 445168 3448 445174 3460
rect 458082 3448 458088 3460
rect 445168 3420 458088 3448
rect 445168 3408 445174 3420
rect 458082 3408 458088 3420
rect 458140 3408 458146 3460
rect 458818 3408 458824 3460
rect 458876 3448 458882 3460
rect 484026 3448 484032 3460
rect 458876 3420 484032 3448
rect 458876 3408 458882 3420
rect 484026 3408 484032 3420
rect 484084 3408 484090 3460
rect 514110 3408 514116 3460
rect 514168 3448 514174 3460
rect 514754 3448 514760 3460
rect 514168 3420 514760 3448
rect 514168 3408 514174 3420
rect 514754 3408 514760 3420
rect 514812 3408 514818 3460
rect 527910 3408 527916 3460
rect 527968 3448 527974 3460
rect 533706 3448 533712 3460
rect 527968 3420 533712 3448
rect 527968 3408 527974 3420
rect 533706 3408 533712 3420
rect 533764 3408 533770 3460
rect 570598 3408 570604 3460
rect 570656 3448 570662 3460
rect 572714 3448 572720 3460
rect 570656 3420 572720 3448
rect 570656 3408 570662 3420
rect 572714 3408 572720 3420
rect 572772 3408 572778 3460
rect 415544 3352 422294 3380
rect 415544 3340 415550 3352
rect 428458 3340 428464 3392
rect 428516 3380 428522 3392
rect 437750 3380 437756 3392
rect 428516 3352 437756 3380
rect 428516 3340 428522 3352
rect 437750 3340 437756 3352
rect 437808 3340 437814 3392
rect 446398 3340 446404 3392
rect 446456 3380 446462 3392
rect 452102 3380 452108 3392
rect 446456 3352 452108 3380
rect 446456 3340 446462 3352
rect 452102 3340 452108 3352
rect 452160 3340 452166 3392
rect 514018 3340 514024 3392
rect 514076 3380 514082 3392
rect 515950 3380 515956 3392
rect 514076 3352 515956 3380
rect 514076 3340 514082 3352
rect 515950 3340 515956 3352
rect 516008 3340 516014 3392
rect 554038 3340 554044 3392
rect 554096 3380 554102 3392
rect 559742 3380 559748 3392
rect 554096 3352 559748 3380
rect 554096 3340 554102 3352
rect 559742 3340 559748 3352
rect 559800 3340 559806 3392
rect 17034 3272 17040 3324
rect 17092 3312 17098 3324
rect 21358 3312 21364 3324
rect 17092 3284 21364 3312
rect 17092 3272 17098 3284
rect 21358 3272 21364 3284
rect 21416 3272 21422 3324
rect 293494 3272 293500 3324
rect 293552 3312 293558 3324
rect 298094 3312 298100 3324
rect 293552 3284 298100 3312
rect 293552 3272 293558 3284
rect 298094 3272 298100 3284
rect 298152 3272 298158 3324
rect 307754 3272 307760 3324
rect 307812 3312 307818 3324
rect 309042 3312 309048 3324
rect 307812 3284 309048 3312
rect 307812 3272 307818 3284
rect 309042 3272 309048 3284
rect 309100 3272 309106 3324
rect 324314 3272 324320 3324
rect 324372 3312 324378 3324
rect 325602 3312 325608 3324
rect 324372 3284 325608 3312
rect 324372 3272 324378 3284
rect 325602 3272 325608 3284
rect 325660 3272 325666 3324
rect 332686 3272 332692 3324
rect 332744 3312 332750 3324
rect 333882 3312 333888 3324
rect 332744 3284 333888 3312
rect 332744 3272 332750 3284
rect 333882 3272 333888 3284
rect 333940 3272 333946 3324
rect 340874 3272 340880 3324
rect 340932 3312 340938 3324
rect 342162 3312 342168 3324
rect 340932 3284 342168 3312
rect 340932 3272 340938 3284
rect 342162 3272 342168 3284
rect 342220 3272 342226 3324
rect 430850 3272 430856 3324
rect 430908 3312 430914 3324
rect 439314 3312 439320 3324
rect 430908 3284 439320 3312
rect 430908 3272 430914 3284
rect 439314 3272 439320 3284
rect 439372 3272 439378 3324
rect 504358 3272 504364 3324
rect 504416 3312 504422 3324
rect 507670 3312 507676 3324
rect 504416 3284 507676 3312
rect 504416 3272 504422 3284
rect 507670 3272 507676 3284
rect 507728 3272 507734 3324
rect 1670 3204 1676 3256
rect 1728 3244 1734 3256
rect 8938 3244 8944 3256
rect 1728 3216 8944 3244
rect 1728 3204 1734 3216
rect 8938 3204 8944 3216
rect 8996 3204 9002 3256
rect 252370 3204 252376 3256
rect 252428 3244 252434 3256
rect 260098 3244 260104 3256
rect 252428 3216 260104 3244
rect 252428 3204 252434 3216
rect 260098 3204 260104 3216
rect 260156 3204 260162 3256
rect 272426 3204 272432 3256
rect 272484 3244 272490 3256
rect 275278 3244 275284 3256
rect 272484 3216 275284 3244
rect 272484 3204 272490 3216
rect 275278 3204 275284 3216
rect 275336 3204 275342 3256
rect 432046 3204 432052 3256
rect 432104 3244 432110 3256
rect 439498 3244 439504 3256
rect 432104 3216 439504 3244
rect 432104 3204 432110 3216
rect 439498 3204 439504 3216
rect 439556 3204 439562 3256
rect 280706 3136 280712 3188
rect 280764 3176 280770 3188
rect 283190 3176 283196 3188
rect 280764 3148 283196 3176
rect 280764 3136 280770 3148
rect 283190 3136 283196 3148
rect 283248 3136 283254 3188
rect 476758 3136 476764 3188
rect 476816 3176 476822 3188
rect 479334 3176 479340 3188
rect 476816 3148 479340 3176
rect 476816 3136 476822 3148
rect 479334 3136 479340 3148
rect 479392 3136 479398 3188
rect 485038 3136 485044 3188
rect 485096 3176 485102 3188
rect 487614 3176 487620 3188
rect 485096 3148 487620 3176
rect 485096 3136 485102 3148
rect 487614 3136 487620 3148
rect 487672 3136 487678 3188
rect 534718 3136 534724 3188
rect 534776 3176 534782 3188
rect 537202 3176 537208 3188
rect 534776 3148 537208 3176
rect 534776 3136 534782 3148
rect 537202 3136 537208 3148
rect 537260 3136 537266 3188
rect 560938 3136 560944 3188
rect 560996 3176 561002 3188
rect 563238 3176 563244 3188
rect 560996 3148 563244 3176
rect 560996 3136 561002 3148
rect 563238 3136 563244 3148
rect 563296 3136 563302 3188
rect 567838 3136 567844 3188
rect 567896 3176 567902 3188
rect 570322 3176 570328 3188
rect 567896 3148 570328 3176
rect 567896 3136 567902 3148
rect 570322 3136 570328 3148
rect 570380 3136 570386 3188
rect 471238 3068 471244 3120
rect 471296 3108 471302 3120
rect 473446 3108 473452 3120
rect 471296 3080 473452 3108
rect 471296 3068 471302 3080
rect 473446 3068 473452 3080
rect 473504 3068 473510 3120
rect 520918 3068 520924 3120
rect 520976 3108 520982 3120
rect 523034 3108 523040 3120
rect 520976 3080 523040 3108
rect 520976 3068 520982 3080
rect 523034 3068 523040 3080
rect 523092 3068 523098 3120
rect 284478 3000 284484 3052
rect 284536 3040 284542 3052
rect 286594 3040 286600 3052
rect 284536 3012 286600 3040
rect 284536 3000 284542 3012
rect 286594 3000 286600 3012
rect 286652 3000 286658 3052
rect 464338 3000 464344 3052
rect 464396 3040 464402 3052
rect 466270 3040 466276 3052
rect 464396 3012 466276 3040
rect 464396 3000 464402 3012
rect 466270 3000 466276 3012
rect 466328 3000 466334 3052
rect 478230 3000 478236 3052
rect 478288 3040 478294 3052
rect 480530 3040 480536 3052
rect 478288 3012 480536 3040
rect 478288 3000 478294 3012
rect 480530 3000 480536 3012
rect 480588 3000 480594 3052
rect 503070 3000 503076 3052
rect 503128 3040 503134 3052
rect 505370 3040 505376 3052
rect 503128 3012 505376 3040
rect 503128 3000 503134 3012
rect 505370 3000 505376 3012
rect 505428 3000 505434 3052
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 10410 2972 10416 2984
rect 8812 2944 10416 2972
rect 8812 2932 8818 2944
rect 10410 2932 10416 2944
rect 10468 2932 10474 2984
rect 19426 2932 19432 2984
rect 19484 2972 19490 2984
rect 25498 2972 25504 2984
rect 19484 2944 25504 2972
rect 19484 2932 19490 2944
rect 25498 2932 25504 2944
rect 25556 2932 25562 2984
rect 457438 2932 457444 2984
rect 457496 2972 457502 2984
rect 459186 2972 459192 2984
rect 457496 2944 459192 2972
rect 457496 2932 457502 2944
rect 459186 2932 459192 2944
rect 459244 2932 459250 2984
rect 494790 2864 494796 2916
rect 494848 2904 494854 2916
rect 499390 2904 499396 2916
rect 494848 2876 499396 2904
rect 494848 2864 494854 2876
rect 499390 2864 499396 2876
rect 499448 2864 499454 2916
rect 273622 2796 273628 2848
rect 273680 2836 273686 2848
rect 278682 2836 278688 2848
rect 273680 2808 278688 2836
rect 273680 2796 273686 2808
rect 278682 2796 278688 2808
rect 278740 2796 278746 2848
rect 316034 1096 316040 1148
rect 316092 1136 316098 1148
rect 317322 1136 317328 1148
rect 316092 1108 317328 1136
rect 316092 1096 316098 1108
rect 317322 1096 317328 1108
rect 317380 1096 317386 1148
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 348792 700544 348844 700596
rect 357716 700544 357768 700596
rect 332508 700476 332560 700528
rect 358820 700476 358872 700528
rect 300124 700408 300176 700460
rect 357624 700408 357676 700460
rect 283840 700340 283892 700392
rect 357532 700340 357584 700392
rect 217968 700272 218020 700324
rect 235172 700272 235224 700324
rect 267648 700272 267700 700324
rect 357440 700272 357492 700324
rect 374644 700272 374696 700324
rect 397460 700272 397512 700324
rect 431224 700272 431276 700324
rect 462320 700272 462372 700324
rect 462964 700272 463016 700324
rect 559656 700272 559708 700324
rect 105452 699728 105504 699780
rect 108304 699728 108356 699780
rect 428464 699660 428516 699712
rect 429844 699660 429896 699712
rect 387064 696940 387116 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 171784 683136 171836 683188
rect 371884 670692 371936 670744
rect 580172 670692 580224 670744
rect 3516 656888 3568 656940
rect 21364 656888 21416 656940
rect 373264 643084 373316 643136
rect 580172 643084 580224 643136
rect 2780 632068 2832 632120
rect 4804 632068 4856 632120
rect 367744 630640 367796 630692
rect 579988 630640 580040 630692
rect 363604 616836 363656 616888
rect 580172 616836 580224 616888
rect 3332 605820 3384 605872
rect 17224 605820 17276 605872
rect 369124 590656 369176 590708
rect 580172 590656 580224 590708
rect 3332 579640 3384 579692
rect 10324 579640 10376 579692
rect 359464 576852 359516 576904
rect 580172 576852 580224 576904
rect 3148 553664 3200 553716
rect 8944 553664 8996 553716
rect 3332 527144 3384 527196
rect 14464 527144 14516 527196
rect 3332 514768 3384 514820
rect 18604 514768 18656 514820
rect 2872 500964 2924 501016
rect 13084 500964 13136 501016
rect 360844 563048 360896 563100
rect 580172 563048 580224 563100
rect 496084 536800 496136 536852
rect 579896 536800 579948 536852
rect 480904 484372 480956 484424
rect 580172 484372 580224 484424
rect 217324 478864 217376 478916
rect 220084 478864 220136 478916
rect 309140 478252 309192 478304
rect 357716 478252 357768 478304
rect 218060 478184 218112 478236
rect 313372 478184 313424 478236
rect 21364 478116 21416 478168
rect 346492 478116 346544 478168
rect 217508 476756 217560 476808
rect 233332 476756 233384 476808
rect 255412 476756 255464 476808
rect 264980 476756 265032 476808
rect 251180 476688 251232 476740
rect 260840 476688 260892 476740
rect 277584 476688 277636 476740
rect 302240 476688 302292 476740
rect 255228 476620 255280 476672
rect 259460 476620 259512 476672
rect 278780 476620 278832 476672
rect 305000 476620 305052 476672
rect 238760 476552 238812 476604
rect 244280 476552 244332 476604
rect 236000 476484 236052 476536
rect 242900 476484 242952 476536
rect 242992 476484 243044 476536
rect 252560 476552 252612 476604
rect 252652 476552 252704 476604
rect 263600 476552 263652 476604
rect 282920 476552 282972 476604
rect 310520 476552 310572 476604
rect 248420 476484 248472 476536
rect 258264 476484 258316 476536
rect 262312 476484 262364 476536
rect 276020 476484 276072 476536
rect 280160 476484 280212 476536
rect 307760 476484 307812 476536
rect 236092 476416 236144 476468
rect 247040 476416 247092 476468
rect 256792 476416 256844 476468
rect 267924 476416 267976 476468
rect 285680 476416 285732 476468
rect 314660 476416 314712 476468
rect 245752 476348 245804 476400
rect 255320 476348 255372 476400
rect 258080 476348 258132 476400
rect 260104 476348 260156 476400
rect 260932 476348 260984 476400
rect 273260 476348 273312 476400
rect 284300 476348 284352 476400
rect 313280 476348 313332 476400
rect 237288 476280 237340 476332
rect 238852 476280 238904 476332
rect 240140 476280 240192 476332
rect 241520 476212 241572 476264
rect 244280 476212 244332 476264
rect 258172 476280 258224 476332
rect 249892 476212 249944 476264
rect 263692 476212 263744 476264
rect 287060 476280 287112 476332
rect 317420 476280 317472 476332
rect 242808 476144 242860 476196
rect 244924 476144 244976 476196
rect 262128 476144 262180 476196
rect 264244 476144 264296 476196
rect 270500 476212 270552 476264
rect 288440 476212 288492 476264
rect 320180 476212 320232 476264
rect 234620 476076 234672 476128
rect 235908 476076 235960 476128
rect 241428 476076 241480 476128
rect 242992 476076 243044 476128
rect 244280 476076 244332 476128
rect 245660 476076 245712 476128
rect 252468 476076 252520 476128
rect 253940 476076 253992 476128
rect 260748 476076 260800 476128
rect 262864 476076 262916 476128
rect 263508 476076 263560 476128
rect 265624 476076 265676 476128
rect 289820 476144 289872 476196
rect 322940 476144 322992 476196
rect 277860 476076 277912 476128
rect 291200 476076 291252 476128
rect 325792 476076 325844 476128
rect 219072 475328 219124 475380
rect 241612 475328 241664 475380
rect 302240 475328 302292 475380
rect 542360 475328 542412 475380
rect 3332 474716 3384 474768
rect 329840 474716 329892 474768
rect 219164 474036 219216 474088
rect 247132 474036 247184 474088
rect 6920 473968 6972 474020
rect 345112 473968 345164 474020
rect 217692 472676 217744 472728
rect 251272 472676 251324 472728
rect 332600 472676 332652 472728
rect 374644 472676 374696 472728
rect 17224 472608 17276 472660
rect 347780 472608 347832 472660
rect 217784 471316 217836 471368
rect 254032 471316 254084 471368
rect 299480 471316 299532 471368
rect 580264 471316 580316 471368
rect 14464 471248 14516 471300
rect 327080 471248 327132 471300
rect 267832 469888 267884 469940
rect 285772 469888 285824 469940
rect 298100 469888 298152 469940
rect 367744 469888 367796 469940
rect 10324 469820 10376 469872
rect 324320 469820 324372 469872
rect 269212 468528 269264 468580
rect 287152 468528 287204 468580
rect 108304 468460 108356 468512
rect 316040 468460 316092 468512
rect 318800 468460 318852 468512
rect 496084 468460 496136 468512
rect 295340 467168 295392 467220
rect 359464 467168 359516 467220
rect 171784 467100 171836 467152
rect 320180 467100 320232 467152
rect 4804 465672 4856 465724
rect 322940 465672 322992 465724
rect 325700 465672 325752 465724
rect 387064 465672 387116 465724
rect 169760 464312 169812 464364
rect 313372 464312 313424 464364
rect 323032 464312 323084 464364
rect 373264 464312 373316 464364
rect 329932 462952 329984 463004
rect 431224 462952 431276 463004
rect 3332 462340 3384 462392
rect 331312 462340 331364 462392
rect 40040 461592 40092 461644
rect 318892 461592 318944 461644
rect 321560 461592 321612 461644
rect 369124 461592 369176 461644
rect 270776 460232 270828 460284
rect 289912 460232 289964 460284
rect 307760 460232 307812 460284
rect 364340 460232 364392 460284
rect 8944 460164 8996 460216
rect 349160 460164 349212 460216
rect 273168 458872 273220 458924
rect 281816 458872 281868 458924
rect 219256 458804 219308 458856
rect 244372 458804 244424 458856
rect 278688 458804 278740 458856
rect 289176 458804 289228 458856
rect 317420 458804 317472 458856
rect 480904 458804 480956 458856
rect 266452 457512 266504 457564
rect 283012 457512 283064 457564
rect 305368 457512 305420 457564
rect 428464 457512 428516 457564
rect 13084 457444 13136 457496
rect 349528 457444 349580 457496
rect 265072 456084 265124 456136
rect 280252 456084 280304 456136
rect 303160 456084 303212 456136
rect 494060 456084 494112 456136
rect 18604 456016 18656 456068
rect 328920 456016 328972 456068
rect 274456 454792 274508 454844
rect 283288 454792 283340 454844
rect 276020 454724 276072 454776
rect 300860 454724 300912 454776
rect 217876 454656 217928 454708
rect 256056 454656 256108 454708
rect 267556 454656 267608 454708
rect 276112 454656 276164 454708
rect 280068 454656 280120 454708
rect 290648 454656 290700 454708
rect 298744 454656 298796 454708
rect 371884 454656 371936 454708
rect 271788 453432 271840 453484
rect 280344 453432 280396 453484
rect 277308 453364 277360 453416
rect 287704 453364 287756 453416
rect 267648 453296 267700 453348
rect 274640 453296 274692 453348
rect 275192 453296 275244 453348
rect 298192 453296 298244 453348
rect 300952 453296 301004 453348
rect 462964 453296 463016 453348
rect 269028 452004 269080 452056
rect 277492 452004 277544 452056
rect 275928 451936 275980 451988
rect 286232 451936 286284 451988
rect 217600 451868 217652 451920
rect 234712 451868 234764 451920
rect 264888 451868 264940 451920
rect 271880 451868 271932 451920
rect 272248 451868 272300 451920
rect 292580 451868 292632 451920
rect 296720 451868 296772 451920
rect 363604 451868 363656 451920
rect 270408 450644 270460 450696
rect 279240 450644 279292 450696
rect 274088 450576 274140 450628
rect 295432 450576 295484 450628
rect 219348 450508 219400 450560
rect 249800 450508 249852 450560
rect 266268 450508 266320 450560
rect 273352 450508 273404 450560
rect 274548 450508 274600 450560
rect 285128 450508 285180 450560
rect 294696 450508 294748 450560
rect 360844 450508 360896 450560
rect 307208 449624 307260 449676
rect 412640 449624 412692 449676
rect 153200 449556 153252 449608
rect 316040 449556 316092 449608
rect 305000 449488 305052 449540
rect 477500 449488 477552 449540
rect 88340 449420 88392 449472
rect 318248 449420 318300 449472
rect 23480 449352 23532 449404
rect 320456 449352 320508 449404
rect 3424 449284 3476 449336
rect 322664 449284 322716 449336
rect 3516 449216 3568 449268
rect 324872 449216 324924 449268
rect 3608 449148 3660 449200
rect 327080 449148 327132 449200
rect 201500 448060 201552 448112
rect 339592 448060 339644 448112
rect 328552 447992 328604 448044
rect 527180 447992 527232 448044
rect 136640 447924 136692 447976
rect 341800 447924 341852 447976
rect 71780 447856 71832 447908
rect 344008 447856 344060 447908
rect 2872 447788 2924 447840
rect 350632 447788 350684 447840
rect 254584 447040 254636 447092
rect 258632 447040 258684 447092
rect 262864 447040 262916 447092
rect 267464 447040 267516 447092
rect 234620 446972 234672 447024
rect 235540 446972 235592 447024
rect 238760 446972 238812 447024
rect 239220 446972 239272 447024
rect 241520 446972 241572 447024
rect 242164 446972 242216 447024
rect 244280 446972 244332 447024
rect 245108 446972 245160 447024
rect 251824 446972 251876 447024
rect 252744 446972 252796 447024
rect 253940 446972 253992 447024
rect 254676 446972 254728 447024
rect 261484 446972 261536 447024
rect 265992 446972 266044 447024
rect 270408 447040 270460 447092
rect 260104 446904 260156 446956
rect 264520 446904 264572 446956
rect 265624 446904 265676 446956
rect 276020 446972 276072 447024
rect 276756 446972 276808 447024
rect 280160 446972 280212 447024
rect 281172 446972 281224 447024
rect 264244 446836 264296 446888
rect 268936 446904 268988 446956
rect 217968 446700 218020 446752
rect 312360 446700 312412 446752
rect 335176 446632 335228 446684
rect 358820 446632 358872 446684
rect 302056 446564 302108 446616
rect 333980 446564 334032 446616
rect 337384 446564 337436 446616
rect 357440 446564 357492 446616
rect 253204 446496 253256 446548
rect 257160 446496 257212 446548
rect 257988 446496 258040 446548
rect 263048 446496 263100 446548
rect 311624 446496 311676 446548
rect 357532 446496 357584 446548
rect 220084 446428 220136 446480
rect 234344 446428 234396 446480
rect 256608 446428 256660 446480
rect 261576 446428 261628 446480
rect 310152 446428 310204 446480
rect 357624 446428 357676 446480
rect 310888 446360 310940 446412
rect 362224 446360 362276 446412
rect 306472 446292 306524 446344
rect 363604 446292 363656 446344
rect 244924 446224 244976 446276
rect 246856 446224 246908 446276
rect 304264 446224 304316 446276
rect 360844 446224 360896 446276
rect 293224 446156 293276 446208
rect 359464 446156 359516 446208
rect 292488 446088 292540 446140
rect 373264 446088 373316 446140
rect 251088 446020 251140 446072
rect 342536 446020 342588 446072
rect 230940 445952 230992 446004
rect 335912 445952 335964 446004
rect 229744 445884 229796 445936
rect 344744 445884 344796 445936
rect 293960 445816 294012 445868
rect 454684 445816 454736 445868
rect 10324 445748 10376 445800
rect 346952 445748 347004 445800
rect 228456 445136 228508 445188
rect 336648 445136 336700 445188
rect 229928 445068 229980 445120
rect 334440 445068 334492 445120
rect 318800 445000 318852 445052
rect 319444 445000 319496 445052
rect 333980 445000 334032 445052
rect 580264 445000 580316 445052
rect 225604 444932 225656 444984
rect 338856 444932 338908 444984
rect 230020 444864 230072 444916
rect 351368 444864 351420 444916
rect 224224 444796 224276 444848
rect 352840 444796 352892 444848
rect 295432 444728 295484 444780
rect 494704 444728 494756 444780
rect 95976 444660 96028 444712
rect 341064 444660 341116 444712
rect 93124 444592 93176 444644
rect 343272 444592 343324 444644
rect 86224 444524 86276 444576
rect 345480 444524 345532 444576
rect 84844 444456 84896 444508
rect 355048 444456 355100 444508
rect 7564 444388 7616 444440
rect 332232 444388 332284 444440
rect 315304 443708 315356 443760
rect 360936 443708 360988 443760
rect 3516 443640 3568 443692
rect 251088 443640 251140 443692
rect 313096 443640 313148 443692
rect 367744 443640 367796 443692
rect 308680 443572 308732 443624
rect 364984 443572 365036 443624
rect 228548 443504 228600 443556
rect 333704 443504 333756 443556
rect 228364 443436 228416 443488
rect 338212 443436 338264 443488
rect 229836 443368 229888 443420
rect 351920 443368 351972 443420
rect 300124 443300 300176 443352
rect 442264 443300 442316 443352
rect 157984 443232 158036 443284
rect 340052 443232 340104 443284
rect 97264 443164 97316 443216
rect 353300 443164 353352 443216
rect 95884 443096 95936 443148
rect 355508 443096 355560 443148
rect 94504 443028 94556 443080
rect 354036 443028 354088 443080
rect 14464 442960 14516 443012
rect 356980 442960 357032 443012
rect 3424 442212 3476 442264
rect 230848 442212 230900 442264
rect 359464 442212 359516 442264
rect 581000 442212 581052 442264
rect 3608 440852 3660 440904
rect 230940 440852 230992 440904
rect 454684 438132 454736 438184
rect 582380 438132 582432 438184
rect 360936 431876 360988 431928
rect 580172 431876 580224 431928
rect 3332 423580 3384 423632
rect 7564 423580 7616 423632
rect 3332 411204 3384 411256
rect 228548 411204 228600 411256
rect 3332 398760 3384 398812
rect 230020 398760 230072 398812
rect 367744 379448 367796 379500
rect 580172 379448 580224 379500
rect 3056 372512 3108 372564
rect 229928 372512 229980 372564
rect 3332 346332 3384 346384
rect 229836 346332 229888 346384
rect 362224 325592 362276 325644
rect 579896 325592 579948 325644
rect 3332 320084 3384 320136
rect 228456 320084 228508 320136
rect 305368 309136 305420 309188
rect 306196 309136 306248 309188
rect 309140 309136 309192 309188
rect 309416 309136 309468 309188
rect 39304 309068 39356 309120
rect 244464 309068 244516 309120
rect 280068 309068 280120 309120
rect 287612 309068 287664 309120
rect 294972 309068 295024 309120
rect 335820 309068 335872 309120
rect 336004 309068 336056 309120
rect 342352 309068 342404 309120
rect 238024 309000 238076 309052
rect 258264 309000 258316 309052
rect 266452 309000 266504 309052
rect 267464 309000 267516 309052
rect 282644 309000 282696 309052
rect 331864 309000 331916 309052
rect 331956 309000 332008 309052
rect 349896 309000 349948 309052
rect 238208 308932 238260 308984
rect 341800 308932 341852 308984
rect 68284 308864 68336 308916
rect 243176 308864 243228 308916
rect 257988 308864 258040 308916
rect 266452 308864 266504 308916
rect 267096 308864 267148 308916
rect 350632 308932 350684 308984
rect 345848 308864 345900 308916
rect 350172 308864 350224 308916
rect 57244 308796 57296 308848
rect 246672 308796 246724 308848
rect 248144 308796 248196 308848
rect 256056 308796 256108 308848
rect 256148 308796 256200 308848
rect 267280 308796 267332 308848
rect 285036 308796 285088 308848
rect 336004 308796 336056 308848
rect 50344 308728 50396 308780
rect 245568 308728 245620 308780
rect 248420 308728 248472 308780
rect 254952 308728 255004 308780
rect 287612 308728 287664 308780
rect 341064 308796 341116 308848
rect 345296 308796 345348 308848
rect 436836 308796 436888 308848
rect 346400 308728 346452 308780
rect 43444 308660 43496 308712
rect 241704 308660 241756 308712
rect 248052 308660 248104 308712
rect 255504 308660 255556 308712
rect 257436 308660 257488 308712
rect 263968 308660 264020 308712
rect 284116 308660 284168 308712
rect 347136 308660 347188 308712
rect 348056 308728 348108 308780
rect 440608 308728 440660 308780
rect 439596 308660 439648 308712
rect 32404 308592 32456 308644
rect 243728 308592 243780 308644
rect 246672 308592 246724 308644
rect 253848 308592 253900 308644
rect 274548 308592 274600 308644
rect 339960 308592 340012 308644
rect 344100 308592 344152 308644
rect 344928 308592 344980 308644
rect 346492 308592 346544 308644
rect 346952 308592 347004 308644
rect 349252 308592 349304 308644
rect 349528 308592 349580 308644
rect 350172 308592 350224 308644
rect 438124 308592 438176 308644
rect 244924 308524 244976 308576
rect 247040 308524 247092 308576
rect 25504 308456 25556 308508
rect 242992 308456 243044 308508
rect 246580 308456 246632 308508
rect 247224 308456 247276 308508
rect 247592 308456 247644 308508
rect 247776 308456 247828 308508
rect 7564 308388 7616 308440
rect 240784 308388 240836 308440
rect 243084 308388 243136 308440
rect 243544 308388 243596 308440
rect 246304 308388 246356 308440
rect 242992 308320 243044 308372
rect 244096 308320 244148 308372
rect 241612 308252 241664 308304
rect 241796 308252 241848 308304
rect 241980 308252 242032 308304
rect 242440 308252 242492 308304
rect 244556 308252 244608 308304
rect 245384 308252 245436 308304
rect 245936 308252 245988 308304
rect 247224 308252 247276 308304
rect 244464 308184 244516 308236
rect 245200 308184 245252 308236
rect 245844 308184 245896 308236
rect 246856 308184 246908 308236
rect 247408 308184 247460 308236
rect 247960 308252 248012 308304
rect 248328 308524 248380 308576
rect 248420 308456 248472 308508
rect 248328 308388 248380 308440
rect 257160 308524 257212 308576
rect 277124 308524 277176 308576
rect 339408 308524 339460 308576
rect 344192 308524 344244 308576
rect 438032 308524 438084 308576
rect 248788 308456 248840 308508
rect 249064 308456 249116 308508
rect 267832 308456 267884 308508
rect 268200 308456 268252 308508
rect 270500 308456 270552 308508
rect 271512 308456 271564 308508
rect 277308 308456 277360 308508
rect 336004 308456 336056 308508
rect 342352 308456 342404 308508
rect 343272 308456 343324 308508
rect 344744 308456 344796 308508
rect 439504 308456 439556 308508
rect 250260 308388 250312 308440
rect 250904 308388 250956 308440
rect 251180 308388 251232 308440
rect 251824 308388 251876 308440
rect 252652 308388 252704 308440
rect 252928 308388 252980 308440
rect 264612 308388 264664 308440
rect 265072 308388 265124 308440
rect 265164 308388 265216 308440
rect 265440 308388 265492 308440
rect 266452 308388 266504 308440
rect 266912 308388 266964 308440
rect 267740 308388 267792 308440
rect 268752 308388 268804 308440
rect 269304 308388 269356 308440
rect 269856 308388 269908 308440
rect 271236 308388 271288 308440
rect 271880 308388 271932 308440
rect 272156 308388 272208 308440
rect 272984 308388 273036 308440
rect 302332 308388 302384 308440
rect 302608 308388 302660 308440
rect 302700 308388 302752 308440
rect 302976 308388 303028 308440
rect 303804 308388 303856 308440
rect 304816 308388 304868 308440
rect 305276 308388 305328 308440
rect 306104 308388 306156 308440
rect 306196 308388 306248 308440
rect 438860 308388 438912 308440
rect 248420 308320 248472 308372
rect 249616 308320 249668 308372
rect 252836 308320 252888 308372
rect 253480 308320 253532 308372
rect 270684 308320 270736 308372
rect 271328 308320 271380 308372
rect 271972 308320 272024 308372
rect 273168 308320 273220 308372
rect 282828 308320 282880 308372
rect 330944 308320 330996 308372
rect 332508 308320 332560 308372
rect 248604 308252 248656 308304
rect 249248 308252 249300 308304
rect 251456 308252 251508 308304
rect 252192 308252 252244 308304
rect 252560 308252 252612 308304
rect 253112 308252 253164 308304
rect 263600 308252 263652 308304
rect 263968 308252 264020 308304
rect 265072 308252 265124 308304
rect 265992 308252 266044 308304
rect 266360 308252 266412 308304
rect 266912 308252 266964 308304
rect 267924 308252 267976 308304
rect 268292 308252 268344 308304
rect 269120 308252 269172 308304
rect 269580 308252 269632 308304
rect 272248 308252 272300 308304
rect 272432 308252 272484 308304
rect 305000 308252 305052 308304
rect 305552 308252 305604 308304
rect 306564 308252 306616 308304
rect 307208 308252 307260 308304
rect 308220 308252 308272 308304
rect 308680 308252 308732 308304
rect 309140 308252 309192 308304
rect 309968 308252 310020 308304
rect 310704 308252 310756 308304
rect 311716 308252 311768 308304
rect 342536 308252 342588 308304
rect 343088 308252 343140 308304
rect 241796 308116 241848 308168
rect 242808 308116 242860 308168
rect 245660 308116 245712 308168
rect 246212 308116 246264 308168
rect 247316 308116 247368 308168
rect 248236 308116 248288 308168
rect 243636 308048 243688 308100
rect 252928 308184 252980 308236
rect 253664 308184 253716 308236
rect 263784 308184 263836 308236
rect 264704 308184 264756 308236
rect 268384 308184 268436 308236
rect 272800 308184 272852 308236
rect 265440 308116 265492 308168
rect 266176 308116 266228 308168
rect 266636 308116 266688 308168
rect 267004 308116 267056 308168
rect 267924 308116 267976 308168
rect 268568 308116 268620 308168
rect 269396 308116 269448 308168
rect 269948 308116 270000 308168
rect 272248 308116 272300 308168
rect 272616 308116 272668 308168
rect 250168 308048 250220 308100
rect 253204 308048 253256 308100
rect 258632 308048 258684 308100
rect 266544 308048 266596 308100
rect 267648 308048 267700 308100
rect 286048 308048 286100 308100
rect 291844 308048 291896 308100
rect 291936 308048 291988 308100
rect 293500 308048 293552 308100
rect 240508 307980 240560 308032
rect 241336 307980 241388 308032
rect 243728 307980 243780 308032
rect 245016 307980 245068 308032
rect 248880 307980 248932 308032
rect 249432 307980 249484 308032
rect 249800 307980 249852 308032
rect 249892 307980 249944 308032
rect 250536 307980 250588 308032
rect 265256 307980 265308 308032
rect 265808 307980 265860 308032
rect 269396 307980 269448 308032
rect 270224 307980 270276 308032
rect 242164 307912 242216 307964
rect 248328 307912 248380 307964
rect 250168 307912 250220 307964
rect 250720 307912 250772 307964
rect 254676 307844 254728 307896
rect 258448 307844 258500 307896
rect 246304 307776 246356 307828
rect 246672 307776 246724 307828
rect 247684 307776 247736 307828
rect 248144 307776 248196 307828
rect 255964 307776 256016 307828
rect 256976 307776 257028 307828
rect 260196 307776 260248 307828
rect 262312 307776 262364 307828
rect 265624 307776 265676 307828
rect 269212 307776 269264 307828
rect 269764 307776 269816 307828
rect 280712 307980 280764 308032
rect 290740 307980 290792 308032
rect 305092 308116 305144 308168
rect 305920 308116 305972 308168
rect 306656 308116 306708 308168
rect 307024 308116 307076 308168
rect 308036 308116 308088 308168
rect 308404 308116 308456 308168
rect 309324 308116 309376 308168
rect 310336 308116 310388 308168
rect 306380 308048 306432 308100
rect 307576 308048 307628 308100
rect 307852 308048 307904 308100
rect 309048 308048 309100 308100
rect 304080 307980 304132 308032
rect 304632 307980 304684 308032
rect 307760 307980 307812 308032
rect 308864 307980 308916 308032
rect 310612 307980 310664 308032
rect 311072 307980 311124 308032
rect 311716 307980 311768 308032
rect 312452 307980 312504 308032
rect 286232 307912 286284 307964
rect 293316 307912 293368 307964
rect 295432 307912 295484 307964
rect 297272 307912 297324 307964
rect 302792 307912 302844 307964
rect 303528 307912 303580 307964
rect 303896 307912 303948 307964
rect 304448 307912 304500 307964
rect 310704 307912 310756 307964
rect 311440 307912 311492 307964
rect 278228 307844 278280 307896
rect 279792 307844 279844 307896
rect 279884 307844 279936 307896
rect 281264 307844 281316 307896
rect 285128 307844 285180 307896
rect 287796 307844 287848 307896
rect 294696 307844 294748 307896
rect 296260 307844 296312 307896
rect 302608 307844 302660 307896
rect 303344 307844 303396 307896
rect 303712 307844 303764 307896
rect 304264 307844 304316 307896
rect 310796 307844 310848 307896
rect 311808 307844 311860 307896
rect 321468 308184 321520 308236
rect 321836 308184 321888 308236
rect 335820 308184 335872 308236
rect 343456 308184 343508 308236
rect 341432 308116 341484 308168
rect 342168 308116 342220 308168
rect 345204 308320 345256 308372
rect 345664 308320 345716 308372
rect 346952 308320 347004 308372
rect 347688 308320 347740 308372
rect 348056 308320 348108 308372
rect 348424 308320 348476 308372
rect 349160 308320 349212 308372
rect 349620 308320 349672 308372
rect 345112 308252 345164 308304
rect 346216 308252 346268 308304
rect 346676 308252 346728 308304
rect 347504 308252 347556 308304
rect 348240 308252 348292 308304
rect 348792 308252 348844 308304
rect 349344 308252 349396 308304
rect 349712 308252 349764 308304
rect 349436 308184 349488 308236
rect 350264 308184 350316 308236
rect 350448 308116 350500 308168
rect 341248 308048 341300 308100
rect 341984 308048 342036 308100
rect 316868 307912 316920 307964
rect 343640 307912 343692 307964
rect 331128 307844 331180 307896
rect 273996 307776 274048 307828
rect 275008 307776 275060 307828
rect 275468 307776 275520 307828
rect 276112 307776 276164 307828
rect 279700 307776 279752 307828
rect 280344 307776 280396 307828
rect 280988 307776 281040 307828
rect 282736 307776 282788 307828
rect 284208 307776 284260 307828
rect 284484 307776 284536 307828
rect 285312 307776 285364 307828
rect 286324 307776 286376 307828
rect 288808 307776 288860 307828
rect 291936 307776 291988 307828
rect 293592 307776 293644 307828
rect 294604 307776 294656 307828
rect 295248 307776 295300 307828
rect 296076 307776 296128 307828
rect 302424 307776 302476 307828
rect 303160 307776 303212 307828
rect 310520 307776 310572 307828
rect 311624 307776 311676 307828
rect 312912 307776 312964 307828
rect 315304 307776 315356 307828
rect 336004 307776 336056 307828
rect 344376 307776 344428 307828
rect 269212 307640 269264 307692
rect 270408 307640 270460 307692
rect 270592 307368 270644 307420
rect 270960 307368 271012 307420
rect 64880 307232 64932 307284
rect 249800 307232 249852 307284
rect 52460 307164 52512 307216
rect 247960 307164 248012 307216
rect 31024 307096 31076 307148
rect 244740 307096 244792 307148
rect 314752 307096 314804 307148
rect 478144 307096 478196 307148
rect 8944 307028 8996 307080
rect 240140 307028 240192 307080
rect 316224 307028 316276 307080
rect 489920 307028 489972 307080
rect 253940 306960 253992 307012
rect 254216 306960 254268 307012
rect 251548 306824 251600 306876
rect 252376 306824 252428 306876
rect 277768 306960 277820 307012
rect 319076 306824 319128 306876
rect 319352 306824 319404 306876
rect 270960 306756 271012 306808
rect 271696 306756 271748 306808
rect 277676 306756 277728 306808
rect 299848 306688 299900 306740
rect 258816 306552 258868 306604
rect 268108 306552 268160 306604
rect 268936 306552 268988 306604
rect 296720 306552 296772 306604
rect 297180 306552 297232 306604
rect 255504 306348 255556 306400
rect 255872 306348 255924 306400
rect 258264 306348 258316 306400
rect 277584 306484 277636 306536
rect 277860 306484 277912 306536
rect 285680 306484 285732 306536
rect 286048 306484 286100 306536
rect 286140 306484 286192 306536
rect 286600 306484 286652 306536
rect 289820 306484 289872 306536
rect 291016 306484 291068 306536
rect 292948 306484 293000 306536
rect 293224 306484 293276 306536
rect 329380 306552 329432 306604
rect 332968 306552 333020 306604
rect 314752 306484 314804 306536
rect 315672 306484 315724 306536
rect 317512 306484 317564 306536
rect 317972 306484 318024 306536
rect 328460 306484 328512 306536
rect 329472 306484 329524 306536
rect 259552 306416 259604 306468
rect 259920 306416 259972 306468
rect 277492 306416 277544 306468
rect 278136 306416 278188 306468
rect 278964 306416 279016 306468
rect 279240 306416 279292 306468
rect 286416 306416 286468 306468
rect 289912 306416 289964 306468
rect 290372 306416 290424 306468
rect 291200 306416 291252 306468
rect 291476 306416 291528 306468
rect 292672 306416 292724 306468
rect 293408 306416 293460 306468
rect 293960 306416 294012 306468
rect 295892 306416 295944 306468
rect 298192 306416 298244 306468
rect 298468 306416 298520 306468
rect 299848 306416 299900 306468
rect 300860 306416 300912 306468
rect 302056 306416 302108 306468
rect 314844 306416 314896 306468
rect 315488 306416 315540 306468
rect 316224 306416 316276 306468
rect 316592 306416 316644 306468
rect 320272 306416 320324 306468
rect 320732 306416 320784 306468
rect 321744 306416 321796 306468
rect 322204 306416 322256 306468
rect 324504 306416 324556 306468
rect 325148 306416 325200 306468
rect 325884 306416 325936 306468
rect 326344 306416 326396 306468
rect 327448 306416 327500 306468
rect 328092 306416 328144 306468
rect 328552 306416 328604 306468
rect 329012 306416 329064 306468
rect 332692 306416 332744 306468
rect 333704 306416 333756 306468
rect 334348 306416 334400 306468
rect 334624 306416 334676 306468
rect 348608 306416 348660 306468
rect 259460 306348 259512 306400
rect 260472 306348 260524 306400
rect 261116 306348 261168 306400
rect 261944 306348 261996 306400
rect 262312 306348 262364 306400
rect 263048 306348 263100 306400
rect 273260 306348 273312 306400
rect 274272 306348 274324 306400
rect 274732 306348 274784 306400
rect 275928 306348 275980 306400
rect 276204 306348 276256 306400
rect 277216 306348 277268 306400
rect 281724 306348 281776 306400
rect 282368 306348 282420 306400
rect 284668 306348 284720 306400
rect 285496 306348 285548 306400
rect 285680 306348 285732 306400
rect 285956 306348 286008 306400
rect 286784 306348 286836 306400
rect 287060 306348 287112 306400
rect 287888 306348 287940 306400
rect 288716 306348 288768 306400
rect 289544 306348 289596 306400
rect 290188 306348 290240 306400
rect 290832 306348 290884 306400
rect 292580 306348 292632 306400
rect 293040 306348 293092 306400
rect 294052 306348 294104 306400
rect 294328 306348 294380 306400
rect 295340 306348 295392 306400
rect 295984 306348 296036 306400
rect 298100 306348 298152 306400
rect 298560 306348 298612 306400
rect 301044 306348 301096 306400
rect 301504 306348 301556 306400
rect 311900 306348 311952 306400
rect 312176 306348 312228 306400
rect 313372 306348 313424 306400
rect 314016 306348 314068 306400
rect 314660 306348 314712 306400
rect 315120 306348 315172 306400
rect 317512 306348 317564 306400
rect 318248 306348 318300 306400
rect 318892 306348 318944 306400
rect 319536 306348 319588 306400
rect 320180 306348 320232 306400
rect 321008 306348 321060 306400
rect 321560 306348 321612 306400
rect 321928 306348 321980 306400
rect 326068 306348 326120 306400
rect 326528 306348 326580 306400
rect 327172 306348 327224 306400
rect 327816 306348 327868 306400
rect 328828 306348 328880 306400
rect 329104 306348 329156 306400
rect 331496 306348 331548 306400
rect 332416 306348 332468 306400
rect 341064 306348 341116 306400
rect 341340 306348 341392 306400
rect 347964 306348 348016 306400
rect 3332 306280 3384 306332
rect 228364 306280 228416 306332
rect 255412 306280 255464 306332
rect 256424 306280 256476 306332
rect 259828 306280 259880 306332
rect 260656 306280 260708 306332
rect 260932 306280 260984 306332
rect 261576 306280 261628 306332
rect 262588 306280 262640 306332
rect 262864 306280 262916 306332
rect 273352 306280 273404 306332
rect 274088 306280 274140 306332
rect 274824 306280 274876 306332
rect 275744 306280 275796 306332
rect 276112 306280 276164 306332
rect 276664 306280 276716 306332
rect 277584 306280 277636 306332
rect 278688 306280 278740 306332
rect 280344 306280 280396 306332
rect 281080 306280 281132 306332
rect 281908 306280 281960 306332
rect 282184 306280 282236 306332
rect 282276 306280 282328 306332
rect 334808 306280 334860 306332
rect 254216 306212 254268 306264
rect 254768 306212 254820 306264
rect 256792 306212 256844 306264
rect 257528 306212 257580 306264
rect 258172 306212 258224 306264
rect 259368 306212 259420 306264
rect 259644 306212 259696 306264
rect 260012 306212 260064 306264
rect 260840 306212 260892 306264
rect 261300 306212 261352 306264
rect 262496 306212 262548 306264
rect 263416 306212 263468 306264
rect 271788 306212 271840 306264
rect 329380 306212 329432 306264
rect 334164 306212 334216 306264
rect 335176 306212 335228 306264
rect 335360 306212 335412 306264
rect 335820 306212 335872 306264
rect 336924 306212 336976 306264
rect 337568 306212 337620 306264
rect 338304 306212 338356 306264
rect 339224 306212 339276 306264
rect 339684 306212 339736 306264
rect 340512 306212 340564 306264
rect 256884 306144 256936 306196
rect 257896 306144 257948 306196
rect 275008 306144 275060 306196
rect 275560 306144 275612 306196
rect 276480 306144 276532 306196
rect 277032 306144 277084 306196
rect 280528 306144 280580 306196
rect 281448 306144 281500 306196
rect 281540 306144 281592 306196
rect 255320 306076 255372 306128
rect 255872 306076 255924 306128
rect 257160 306076 257212 306128
rect 257712 306076 257764 306128
rect 259644 306076 259696 306128
rect 260288 306076 260340 306128
rect 260840 306076 260892 306128
rect 262128 306076 262180 306128
rect 271696 306076 271748 306128
rect 332232 306076 332284 306128
rect 335544 306076 335596 306128
rect 273628 306008 273680 306060
rect 274456 306008 274508 306060
rect 276296 306008 276348 306060
rect 276848 306008 276900 306060
rect 277768 306008 277820 306060
rect 278504 306008 278556 306060
rect 278596 306008 278648 306060
rect 344560 306008 344612 306060
rect 255596 305940 255648 305992
rect 256608 305940 256660 305992
rect 256976 305940 257028 305992
rect 257344 305940 257396 305992
rect 275284 305940 275336 305992
rect 345020 305940 345072 305992
rect 255688 305872 255740 305924
rect 256240 305872 256292 305924
rect 272616 305872 272668 305924
rect 345112 305872 345164 305924
rect 272524 305804 272576 305856
rect 345204 305804 345256 305856
rect 88984 305736 89036 305788
rect 253296 305736 253348 305788
rect 269856 305736 269908 305788
rect 347320 305736 347372 305788
rect 71780 305668 71832 305720
rect 251272 305668 251324 305720
rect 270040 305668 270092 305720
rect 347780 305668 347832 305720
rect 35164 305600 35216 305652
rect 244464 305600 244516 305652
rect 267004 305600 267056 305652
rect 347872 305600 347924 305652
rect 257344 305532 257396 305584
rect 257988 305532 258040 305584
rect 275376 305532 275428 305584
rect 278596 305532 278648 305584
rect 279424 305532 279476 305584
rect 279884 305532 279936 305584
rect 281448 305532 281500 305584
rect 274548 305464 274600 305516
rect 281540 305464 281592 305516
rect 284576 305464 284628 305516
rect 284944 305464 284996 305516
rect 285864 305464 285916 305516
rect 286968 305464 287020 305516
rect 287152 305464 287204 305516
rect 287520 305464 287572 305516
rect 288440 305464 288492 305516
rect 288900 305464 288952 305516
rect 290096 305464 290148 305516
rect 290648 305464 290700 305516
rect 291384 305464 291436 305516
rect 291752 305464 291804 305516
rect 292396 305464 292448 305516
rect 274364 305396 274416 305448
rect 282276 305396 282328 305448
rect 288624 305396 288676 305448
rect 289728 305396 289780 305448
rect 289912 305396 289964 305448
rect 290464 305396 290516 305448
rect 291568 305396 291620 305448
rect 292120 305396 292172 305448
rect 294052 305396 294104 305448
rect 295064 305396 295116 305448
rect 295524 305396 295576 305448
rect 296168 305396 296220 305448
rect 296996 305396 297048 305448
rect 297640 305396 297692 305448
rect 298376 305396 298428 305448
rect 299296 305396 299348 305448
rect 299664 305396 299716 305448
rect 300032 305396 300084 305448
rect 301228 305396 301280 305448
rect 301872 305396 301924 305448
rect 278044 305328 278096 305380
rect 278228 305328 278280 305380
rect 287152 305328 287204 305380
rect 288072 305328 288124 305380
rect 288440 305328 288492 305380
rect 289176 305328 289228 305380
rect 291292 305328 291344 305380
rect 292304 305328 292356 305380
rect 299572 305328 299624 305380
rect 300584 305328 300636 305380
rect 301136 305328 301188 305380
rect 301688 305328 301740 305380
rect 277952 305260 278004 305312
rect 278320 305260 278372 305312
rect 299480 305260 299532 305312
rect 300400 305260 300452 305312
rect 298284 305192 298336 305244
rect 298744 305192 298796 305244
rect 332048 305396 332100 305448
rect 313648 305328 313700 305380
rect 313832 305328 313884 305380
rect 316040 305328 316092 305380
rect 316408 305328 316460 305380
rect 317788 305328 317840 305380
rect 318616 305328 318668 305380
rect 318984 305328 319036 305380
rect 319260 305328 319312 305380
rect 320548 305328 320600 305380
rect 321376 305328 321428 305380
rect 321836 305328 321888 305380
rect 322296 305328 322348 305380
rect 323308 305328 323360 305380
rect 324136 305328 324188 305380
rect 324320 305328 324372 305380
rect 324596 305328 324648 305380
rect 324872 305328 324924 305380
rect 325608 305328 325660 305380
rect 326160 305328 326212 305380
rect 326712 305328 326764 305380
rect 327080 305328 327132 305380
rect 327632 305328 327684 305380
rect 328736 305328 328788 305380
rect 329656 305328 329708 305380
rect 332416 305532 332468 305584
rect 337200 305532 337252 305584
rect 336280 305396 336332 305448
rect 333888 305328 333940 305380
rect 316316 305260 316368 305312
rect 317144 305260 317196 305312
rect 318800 305260 318852 305312
rect 319168 305260 319220 305312
rect 320364 305260 320416 305312
rect 321192 305260 321244 305312
rect 321652 305260 321704 305312
rect 322480 305260 322532 305312
rect 322940 305260 322992 305312
rect 323492 305260 323544 305312
rect 325792 305260 325844 305312
rect 326896 305260 326948 305312
rect 327264 305260 327316 305312
rect 328368 305260 328420 305312
rect 328552 305260 328604 305312
rect 329288 305260 329340 305312
rect 296536 305124 296588 305176
rect 316408 305192 316460 305244
rect 317328 305192 317380 305244
rect 318984 305192 319036 305244
rect 319904 305192 319956 305244
rect 321744 305192 321796 305244
rect 322848 305192 322900 305244
rect 323216 305192 323268 305244
rect 323952 305192 324004 305244
rect 324596 305192 324648 305244
rect 325424 305192 325476 305244
rect 327080 305192 327132 305244
rect 328184 305192 328236 305244
rect 299940 305124 299992 305176
rect 300768 305124 300820 305176
rect 318800 305124 318852 305176
rect 320088 305124 320140 305176
rect 322112 305124 322164 305176
rect 322664 305124 322716 305176
rect 322940 305124 322992 305176
rect 323768 305124 323820 305176
rect 282920 305056 282972 305108
rect 284024 305056 284076 305108
rect 294144 305056 294196 305108
rect 294512 305056 294564 305108
rect 296812 304920 296864 304972
rect 297456 304920 297508 304972
rect 278872 304648 278924 304700
rect 279976 304648 280028 304700
rect 313556 304580 313608 304632
rect 314200 304580 314252 304632
rect 313464 304512 313516 304564
rect 314384 304512 314436 304564
rect 91100 304376 91152 304428
rect 253940 304376 253992 304428
rect 317420 304376 317472 304428
rect 318432 304376 318484 304428
rect 18604 304308 18656 304360
rect 241612 304308 241664 304360
rect 254400 304308 254452 304360
rect 254584 304308 254636 304360
rect 315856 304308 315908 304360
rect 485044 304308 485096 304360
rect 13084 304240 13136 304292
rect 240232 304240 240284 304292
rect 254124 304240 254176 304292
rect 255136 304240 255188 304292
rect 292488 304240 292540 304292
rect 292948 304240 293000 304292
rect 319352 304240 319404 304292
rect 507860 304240 507912 304292
rect 335636 303832 335688 303884
rect 336648 303832 336700 303884
rect 312176 303764 312228 303816
rect 312544 303764 312596 303816
rect 311992 303696 312044 303748
rect 312728 303696 312780 303748
rect 312084 303628 312136 303680
rect 313096 303628 313148 303680
rect 282644 303560 282696 303612
rect 330760 303560 330812 303612
rect 271604 303492 271656 303544
rect 337752 303492 337804 303544
rect 261668 303424 261720 303476
rect 334992 303424 335044 303476
rect 258908 303356 258960 303408
rect 335544 303356 335596 303408
rect 258816 303288 258868 303340
rect 336464 303288 336516 303340
rect 338396 303288 338448 303340
rect 338672 303288 338724 303340
rect 258724 303220 258776 303272
rect 337292 303220 337344 303272
rect 256148 303152 256200 303204
rect 337936 303152 337988 303204
rect 267188 303084 267240 303136
rect 348976 303084 349028 303136
rect 82820 303016 82872 303068
rect 252652 303016 252704 303068
rect 256240 303016 256292 303068
rect 338580 303016 338632 303068
rect 27620 302948 27672 303000
rect 244648 302948 244700 303000
rect 264336 302948 264388 303000
rect 349252 302948 349304 303000
rect 17224 302880 17276 302932
rect 241152 302880 241204 302932
rect 261576 302880 261628 302932
rect 350080 302880 350132 302932
rect 286692 302812 286744 302864
rect 332600 302812 332652 302864
rect 283104 302744 283156 302796
rect 283656 302744 283708 302796
rect 285496 302744 285548 302796
rect 331680 302744 331732 302796
rect 293684 302676 293736 302728
rect 331404 302676 331456 302728
rect 338120 302336 338172 302388
rect 338580 302336 338632 302388
rect 294420 302200 294472 302252
rect 294604 302200 294656 302252
rect 308496 301520 308548 301572
rect 440240 301520 440292 301572
rect 39396 301452 39448 301504
rect 245752 301452 245804 301504
rect 317880 301452 317932 301504
rect 500224 301452 500276 301504
rect 289544 300704 289596 300756
rect 334716 300704 334768 300756
rect 288072 300636 288124 300688
rect 333520 300636 333572 300688
rect 286876 300568 286928 300620
rect 333152 300568 333204 300620
rect 285404 300500 285456 300552
rect 331496 300500 331548 300552
rect 284116 300432 284168 300484
rect 341616 300432 341668 300484
rect 279976 300364 280028 300416
rect 338856 300364 338908 300416
rect 277124 300296 277176 300348
rect 339684 300296 339736 300348
rect 310152 300228 310204 300280
rect 449900 300228 449952 300280
rect 71044 300160 71096 300212
rect 249892 300160 249944 300212
rect 317788 300160 317840 300212
rect 502984 300160 503036 300212
rect 21364 300092 21416 300144
rect 242624 300092 242676 300144
rect 327632 300092 327684 300144
rect 554044 300092 554096 300144
rect 70400 298868 70452 298920
rect 251088 298868 251140 298920
rect 53840 298800 53892 298852
rect 248512 298800 248564 298852
rect 312360 298800 312412 298852
rect 462964 298800 463016 298852
rect 22744 298732 22796 298784
rect 243176 298732 243228 298784
rect 319352 298732 319404 298784
rect 512000 298732 512052 298784
rect 238300 297576 238352 297628
rect 342904 297576 342956 297628
rect 92480 297508 92532 297560
rect 254492 297508 254544 297560
rect 57980 297440 58032 297492
rect 248788 297440 248840 297492
rect 35900 297372 35952 297424
rect 246212 297372 246264 297424
rect 320640 297372 320692 297424
rect 516784 297372 516836 297424
rect 80060 296012 80112 296064
rect 253112 296012 253164 296064
rect 320548 296012 320600 296064
rect 520924 296012 520976 296064
rect 60740 295944 60792 295996
rect 248420 295944 248472 295996
rect 329012 295944 329064 295996
rect 566464 295944 566516 295996
rect 310980 294788 311032 294840
rect 453304 294788 453356 294840
rect 319260 294720 319312 294772
rect 504364 294720 504416 294772
rect 69020 294652 69072 294704
rect 250168 294652 250220 294704
rect 323492 294652 323544 294704
rect 527824 294652 527876 294704
rect 12440 294584 12492 294636
rect 241888 294584 241940 294636
rect 324964 294584 325016 294636
rect 542360 294584 542412 294636
rect 3332 293904 3384 293956
rect 224224 293904 224276 293956
rect 323400 293292 323452 293344
rect 534724 293292 534776 293344
rect 93860 293224 93912 293276
rect 254216 293224 254268 293276
rect 328920 293224 328972 293276
rect 571340 293224 571392 293276
rect 98000 291864 98052 291916
rect 255872 291864 255924 291916
rect 313924 291864 313976 291916
rect 476764 291864 476816 291916
rect 75920 291796 75972 291848
rect 251180 291796 251232 291848
rect 323308 291796 323360 291848
rect 538864 291796 538916 291848
rect 78680 290504 78732 290556
rect 251548 290504 251600 290556
rect 22100 290436 22152 290488
rect 243084 290436 243136 290488
rect 327540 290436 327592 290488
rect 563704 290436 563756 290488
rect 85580 289144 85632 289196
rect 252836 289144 252888 289196
rect 30380 289076 30432 289128
rect 244832 289076 244884 289128
rect 328828 289076 328880 289128
rect 570604 289076 570656 289128
rect 308220 287716 308272 287768
rect 440332 287716 440384 287768
rect 34520 287648 34572 287700
rect 244556 287648 244608 287700
rect 328736 287648 328788 287700
rect 575480 287648 575532 287700
rect 309508 286424 309560 286476
rect 442356 286424 442408 286476
rect 309600 286356 309652 286408
rect 448520 286356 448572 286408
rect 49700 286288 49752 286340
rect 247408 286288 247460 286340
rect 326252 286288 326304 286340
rect 553400 286288 553452 286340
rect 312544 285064 312596 285116
rect 454040 285064 454092 285116
rect 63500 284996 63552 285048
rect 250076 284996 250128 285048
rect 313832 284996 313884 285048
rect 471244 284996 471296 285048
rect 26240 284928 26292 284980
rect 242992 284928 243044 284980
rect 327448 284928 327500 284980
rect 560944 284928 560996 284980
rect 77300 283636 77352 283688
rect 251456 283636 251508 283688
rect 313648 283636 313700 283688
rect 471980 283636 472032 283688
rect 40040 283568 40092 283620
rect 245936 283568 245988 283620
rect 313740 283568 313792 283620
rect 473452 283568 473504 283620
rect 310888 282276 310940 282328
rect 452660 282276 452712 282328
rect 81440 282208 81492 282260
rect 252744 282208 252796 282260
rect 310796 282208 310848 282260
rect 460940 282208 460992 282260
rect 44180 282140 44232 282192
rect 245844 282140 245896 282192
rect 319168 282140 319220 282192
rect 506572 282140 506624 282192
rect 309416 280848 309468 280900
rect 444380 280848 444432 280900
rect 4896 280780 4948 280832
rect 240324 280780 240376 280832
rect 319076 280780 319128 280832
rect 509240 280780 509292 280832
rect 309324 279488 309376 279540
rect 446404 279488 446456 279540
rect 10416 279420 10468 279472
rect 240508 279420 240560 279472
rect 317696 279420 317748 279472
rect 499580 279420 499632 279472
rect 310704 278060 310756 278112
rect 457444 278060 457496 278112
rect 320456 277992 320508 278044
rect 517520 277992 517572 278044
rect 312268 276700 312320 276752
rect 460204 276700 460256 276752
rect 320364 276632 320416 276684
rect 521660 276632 521712 276684
rect 312176 275340 312228 275392
rect 464344 275340 464396 275392
rect 55220 275272 55272 275324
rect 248696 275272 248748 275324
rect 323216 275272 323268 275324
rect 539692 275272 539744 275324
rect 59360 273912 59412 273964
rect 248604 273912 248656 273964
rect 312084 273912 312136 273964
rect 467104 273912 467156 273964
rect 364984 273164 365036 273216
rect 579896 273164 579948 273216
rect 62120 272484 62172 272536
rect 249984 272484 250036 272536
rect 308128 271328 308180 271380
rect 436744 271328 436796 271380
rect 313556 271260 313608 271312
rect 475384 271260 475436 271312
rect 327356 271192 327408 271244
rect 560300 271192 560352 271244
rect 66260 271124 66312 271176
rect 250352 271124 250404 271176
rect 328644 271124 328696 271176
rect 567844 271124 567896 271176
rect 314936 269968 314988 270020
rect 481640 269968 481692 270020
rect 326160 269900 326212 269952
rect 556160 269900 556212 269952
rect 327264 269832 327316 269884
rect 567200 269832 567252 269884
rect 73160 269764 73212 269816
rect 251364 269764 251416 269816
rect 328552 269764 328604 269816
rect 571984 269764 572036 269816
rect 313372 268676 313424 268728
rect 474740 268676 474792 268728
rect 313464 268608 313516 268660
rect 477500 268608 477552 268660
rect 314844 268540 314896 268592
rect 484400 268540 484452 268592
rect 322204 268472 322256 268524
rect 524420 268472 524472 268524
rect 324780 268404 324832 268456
rect 546500 268404 546552 268456
rect 77392 268336 77444 268388
rect 251732 268336 251784 268388
rect 324872 268336 324924 268388
rect 549260 268336 549312 268388
rect 2964 267656 3016 267708
rect 225604 267656 225656 267708
rect 314752 267112 314804 267164
rect 485780 267112 485832 267164
rect 316500 267044 316552 267096
rect 492680 267044 492732 267096
rect 317604 266976 317656 267028
rect 494796 266976 494848 267028
rect 84200 265684 84252 265736
rect 253020 265684 253072 265736
rect 316408 265684 316460 265736
rect 496820 265684 496872 265736
rect 7656 265616 7708 265668
rect 240416 265616 240468 265668
rect 317512 265616 317564 265668
rect 502340 265616 502392 265668
rect 317420 264324 317472 264376
rect 503720 264324 503772 264376
rect 318984 264256 319036 264308
rect 511264 264256 511316 264308
rect 17960 264188 18012 264240
rect 241796 264188 241848 264240
rect 326068 264188 326120 264240
rect 556252 264188 556304 264240
rect 318892 263100 318944 263152
rect 510620 263100 510672 263152
rect 320272 263032 320324 263084
rect 516140 263032 516192 263084
rect 324688 262964 324740 263016
rect 545120 262964 545172 263016
rect 324596 262896 324648 262948
rect 547880 262896 547932 262948
rect 41420 262828 41472 262880
rect 246120 262828 246172 262880
rect 325976 262828 326028 262880
rect 552020 262828 552072 262880
rect 320180 261672 320232 261724
rect 520280 261672 520332 261724
rect 322112 261604 322164 261656
rect 531320 261604 531372 261656
rect 323124 261536 323176 261588
rect 535460 261536 535512 261588
rect 324504 261468 324556 261520
rect 540980 261468 541032 261520
rect 311992 260312 312044 260364
rect 466460 260312 466512 260364
rect 316316 260244 316368 260296
rect 495440 260244 495492 260296
rect 322020 260176 322072 260228
rect 527180 260176 527232 260228
rect 11704 260108 11756 260160
rect 241704 260108 241756 260160
rect 363604 260108 363656 260160
rect 580448 260108 580500 260160
rect 313280 258884 313332 258936
rect 470600 258884 470652 258936
rect 316132 258816 316184 258868
rect 488540 258816 488592 258868
rect 316224 258748 316276 258800
rect 491300 258748 491352 258800
rect 56600 258680 56652 258732
rect 248972 258680 249024 258732
rect 360844 258680 360896 258732
rect 580356 258680 580408 258732
rect 321928 257320 321980 257372
rect 523132 257320 523184 257372
rect 297916 256096 297968 256148
rect 330116 256096 330168 256148
rect 297640 256028 297692 256080
rect 332692 256028 332744 256080
rect 297272 255960 297324 256012
rect 336924 255960 336976 256012
rect 3148 255212 3200 255264
rect 157984 255212 158036 255264
rect 238484 254532 238536 254584
rect 346768 254532 346820 254584
rect 373264 254532 373316 254584
rect 581092 254532 581144 254584
rect 60832 253172 60884 253224
rect 248880 253172 248932 253224
rect 307852 253172 307904 253224
rect 443000 253172 443052 253224
rect 315304 251948 315356 252000
rect 467840 251948 467892 252000
rect 321836 251880 321888 251932
rect 528560 251880 528612 251932
rect 74540 251812 74592 251864
rect 251640 251812 251692 251864
rect 321744 251812 321796 251864
rect 531412 251812 531464 251864
rect 288348 251132 288400 251184
rect 334072 251132 334124 251184
rect 293592 251064 293644 251116
rect 339592 251064 339644 251116
rect 292396 250996 292448 251048
rect 339960 250996 340012 251048
rect 290924 250928 290976 250980
rect 338304 250928 338356 250980
rect 291016 250860 291068 250912
rect 338396 250860 338448 250912
rect 275928 250792 275980 250844
rect 331956 250792 332008 250844
rect 349436 250792 349488 250844
rect 438216 250792 438268 250844
rect 283932 250724 283984 250776
rect 342444 250724 342496 250776
rect 349344 250724 349396 250776
rect 441712 250724 441764 250776
rect 281264 250656 281316 250708
rect 342536 250656 342588 250708
rect 349620 250656 349672 250708
rect 441804 250656 441856 250708
rect 310612 250588 310664 250640
rect 456892 250588 456944 250640
rect 310520 250520 310572 250572
rect 459560 250520 459612 250572
rect 13820 250452 13872 250504
rect 242072 250452 242124 250504
rect 318800 250452 318852 250504
rect 514116 250452 514168 250504
rect 296444 250384 296496 250436
rect 341156 250384 341208 250436
rect 289636 250316 289688 250368
rect 334164 250316 334216 250368
rect 299296 250248 299348 250300
rect 341064 250248 341116 250300
rect 296904 249432 296956 249484
rect 297364 249432 297416 249484
rect 309232 249228 309284 249280
rect 445760 249228 445812 249280
rect 314660 249160 314712 249212
rect 481732 249160 481784 249212
rect 297180 249092 297232 249144
rect 325884 249092 325936 249144
rect 554780 249092 554832 249144
rect 325792 249024 325844 249076
rect 557540 249024 557592 249076
rect 297180 248820 297232 248872
rect 293408 248344 293460 248396
rect 303988 248344 304040 248396
rect 298836 248276 298888 248328
rect 348240 248276 348292 248328
rect 282552 248208 282604 248260
rect 337200 248208 337252 248260
rect 346492 248208 346544 248260
rect 436928 248208 436980 248260
rect 278596 248140 278648 248192
rect 341432 248140 341484 248192
rect 346676 248140 346728 248192
rect 438308 248140 438360 248192
rect 278688 248072 278740 248124
rect 346584 248072 346636 248124
rect 347964 248072 348016 248124
rect 441896 248072 441948 248124
rect 283932 248004 283984 248056
rect 304172 248004 304224 248056
rect 305552 248004 305604 248056
rect 437480 248004 437532 248056
rect 286600 247936 286652 247988
rect 302884 247936 302936 247988
rect 305368 247936 305420 247988
rect 437572 247936 437624 247988
rect 287796 247868 287848 247920
rect 302608 247868 302660 247920
rect 306932 247868 306984 247920
rect 440424 247868 440476 247920
rect 289176 247800 289228 247852
rect 302792 247800 302844 247852
rect 305460 247800 305512 247852
rect 438952 247800 439004 247852
rect 285036 247732 285088 247784
rect 302700 247732 302752 247784
rect 306840 247732 306892 247784
rect 440516 247732 440568 247784
rect 31760 247664 31812 247716
rect 243728 247664 243780 247716
rect 304080 247664 304132 247716
rect 439044 247664 439096 247716
rect 296352 247596 296404 247648
rect 342352 247596 342404 247648
rect 293500 247528 293552 247580
rect 338580 247528 338632 247580
rect 297272 247460 297324 247512
rect 334348 247460 334400 247512
rect 288256 247392 288308 247444
rect 335636 247392 335688 247444
rect 295064 247052 295116 247104
rect 298560 247052 298612 247104
rect 295156 246984 295208 247036
rect 349528 246984 349580 247036
rect 277032 246916 277084 246968
rect 331864 246916 331916 246968
rect 281356 246848 281408 246900
rect 343732 246848 343784 246900
rect 275836 246780 275888 246832
rect 344100 246780 344152 246832
rect 274272 246712 274324 246764
rect 345480 246712 345532 246764
rect 273168 246644 273220 246696
rect 348148 246644 348200 246696
rect 350632 246644 350684 246696
rect 439688 246644 439740 246696
rect 309140 246576 309192 246628
rect 448612 246576 448664 246628
rect 316040 246508 316092 246560
rect 490012 246508 490064 246560
rect 322940 246440 322992 246492
rect 538220 246440 538272 246492
rect 324320 246372 324372 246424
rect 543740 246372 543792 246424
rect 95240 246304 95292 246356
rect 243636 246304 243688 246356
rect 285588 246304 285640 246356
rect 292948 246304 293000 246356
rect 327172 246304 327224 246356
rect 564532 246304 564584 246356
rect 298008 246236 298060 246288
rect 346952 246236 347004 246288
rect 297456 246168 297508 246220
rect 336004 246168 336056 246220
rect 299020 246100 299072 246152
rect 335820 246100 335872 246152
rect 296812 245556 296864 245608
rect 298744 245556 298796 245608
rect 306748 245556 306800 245608
rect 437756 245556 437808 245608
rect 295248 245488 295300 245540
rect 302332 245488 302384 245540
rect 306472 245488 306524 245540
rect 437848 245488 437900 245540
rect 290832 245420 290884 245472
rect 303712 245420 303764 245472
rect 305092 245420 305144 245472
rect 437664 245420 437716 245472
rect 292120 245352 292172 245404
rect 302424 245352 302476 245404
rect 306656 245352 306708 245404
rect 439320 245352 439372 245404
rect 293776 245284 293828 245336
rect 301044 245284 301096 245336
rect 306564 245284 306616 245336
rect 439412 245284 439464 245336
rect 305000 245216 305052 245268
rect 437940 245216 437992 245268
rect 296628 245148 296680 245200
rect 303620 245148 303672 245200
rect 305276 245148 305328 245200
rect 439136 245148 439188 245200
rect 305184 245080 305236 245132
rect 439228 245080 439280 245132
rect 291108 245012 291160 245064
rect 302240 245012 302292 245064
rect 311900 245012 311952 245064
rect 463700 245012 463752 245064
rect 321560 244944 321612 244996
rect 525800 244944 525852 244996
rect 3608 244876 3660 244928
rect 229744 244876 229796 244928
rect 293408 244876 293460 244928
rect 300860 244876 300912 244928
rect 329932 244876 329984 244928
rect 576860 244876 576912 244928
rect 279884 244808 279936 244860
rect 345572 244808 345624 244860
rect 297548 244740 297600 244792
rect 337108 244740 337160 244792
rect 299112 244672 299164 244724
rect 332968 244672 333020 244724
rect 288164 244604 288216 244656
rect 295248 244604 295300 244656
rect 299848 244604 299900 244656
rect 297732 244536 297784 244588
rect 330208 244536 330260 244588
rect 293868 244468 293920 244520
rect 300952 244468 301004 244520
rect 301136 244400 301188 244452
rect 291752 244332 291804 244384
rect 297364 244332 297416 244384
rect 297824 243788 297876 243840
rect 316776 243788 316828 243840
rect 299204 243720 299256 243772
rect 338488 243720 338540 243772
rect 290832 243652 290884 243704
rect 335728 243652 335780 243704
rect 294972 243584 295024 243636
rect 342628 243584 342680 243636
rect 286784 243516 286836 243568
rect 341248 243516 341300 243568
rect 97724 243448 97776 243500
rect 297088 243448 297140 243500
rect 97816 243380 97868 243432
rect 297364 243380 297416 243432
rect 297548 243380 297600 243432
rect 3240 241408 3292 241460
rect 97264 241408 97316 241460
rect 3332 215228 3384 215280
rect 95976 215228 96028 215280
rect 3148 188980 3200 189032
rect 94504 188980 94556 189032
rect 3516 164160 3568 164212
rect 93124 164160 93176 164212
rect 297272 243108 297324 243160
rect 297548 243108 297600 243160
rect 293500 239776 293552 239828
rect 293776 239776 293828 239828
rect 297180 195984 297232 196036
rect 298836 195984 298888 196036
rect 295156 195916 295208 195968
rect 297272 195916 297324 195968
rect 280988 193808 281040 193860
rect 297456 193808 297508 193860
rect 283564 191836 283616 191888
rect 299020 191836 299072 191888
rect 297272 189864 297324 189916
rect 298376 189864 298428 189916
rect 238116 174632 238168 174684
rect 260012 174632 260064 174684
rect 245752 174564 245804 174616
rect 277952 174564 278004 174616
rect 237380 174496 237432 174548
rect 276480 174496 276532 174548
rect 239404 173136 239456 173188
rect 266820 173136 266872 173188
rect 282644 171028 282696 171080
rect 297640 171028 297692 171080
rect 297180 170552 297232 170604
rect 298560 170552 298612 170604
rect 238392 170348 238444 170400
rect 282644 170348 282696 170400
rect 293776 168308 293828 168360
rect 297640 168308 297692 168360
rect 238576 167628 238628 167680
rect 297916 167628 297968 167680
rect 97448 159876 97500 159928
rect 297548 159876 297600 159928
rect 97540 159808 97592 159860
rect 297456 159808 297508 159860
rect 97724 159740 97776 159792
rect 283564 159740 283616 159792
rect 97816 159672 97868 159724
rect 280988 159672 281040 159724
rect 97908 159604 97960 159656
rect 238576 159604 238628 159656
rect 286140 159604 286192 159656
rect 299480 159604 299532 159656
rect 97356 159536 97408 159588
rect 238392 159536 238444 159588
rect 287520 159536 287572 159588
rect 302240 159536 302292 159588
rect 288256 159468 288308 159520
rect 336004 159468 336056 159520
rect 289636 159400 289688 159452
rect 338488 159400 338540 159452
rect 173440 159332 173492 159384
rect 294696 159332 294748 159384
rect 297640 159332 297692 159384
rect 348240 159332 348292 159384
rect 291016 159264 291068 159316
rect 351000 159264 351052 159316
rect 290924 159196 290976 159248
rect 353576 159196 353628 159248
rect 206008 159128 206060 159180
rect 267096 159128 267148 159180
rect 293592 159128 293644 159180
rect 356060 159128 356112 159180
rect 165988 159060 166040 159112
rect 238208 159060 238260 159112
rect 299296 159060 299348 159112
rect 363512 159060 363564 159112
rect 156052 158992 156104 159044
rect 243544 158992 243596 159044
rect 296444 158992 296496 159044
rect 360936 158992 360988 159044
rect 158536 158924 158588 158976
rect 257528 158924 257580 158976
rect 281264 158924 281316 158976
rect 370964 158924 371016 158976
rect 284024 158856 284076 158908
rect 368204 158856 368256 158908
rect 168288 158788 168340 158840
rect 284944 158788 284996 158840
rect 292396 158788 292448 158840
rect 358452 158788 358504 158840
rect 160928 158720 160980 158772
rect 289084 158720 289136 158772
rect 297824 158720 297876 158772
rect 373356 158720 373408 158772
rect 120632 158652 120684 158704
rect 288072 158652 288124 158704
rect 288256 158652 288308 158704
rect 290832 158652 290884 158704
rect 340972 158652 341024 158704
rect 376024 158652 376076 158704
rect 438032 158652 438084 158704
rect 282552 158584 282604 158636
rect 345940 158584 345992 158636
rect 378600 158584 378652 158636
rect 439504 158584 439556 158636
rect 119712 158516 119764 158568
rect 286140 158516 286192 158568
rect 286692 158516 286744 158568
rect 286784 158516 286836 158568
rect 365812 158516 365864 158568
rect 380992 158516 381044 158568
rect 436836 158516 436888 158568
rect 288164 158448 288216 158500
rect 343548 158448 343600 158500
rect 383568 158448 383620 158500
rect 438124 158448 438176 158500
rect 126520 158380 126572 158432
rect 292304 158380 292356 158432
rect 293684 158380 293736 158432
rect 328276 158380 328328 158432
rect 385960 158380 386012 158432
rect 439596 158380 439648 158432
rect 133512 158312 133564 158364
rect 299204 158312 299256 158364
rect 333428 158312 333480 158364
rect 388536 158312 388588 158364
rect 436928 158312 436980 158364
rect 130568 158244 130620 158296
rect 281448 158244 281500 158296
rect 329932 158244 329984 158296
rect 391480 158244 391532 158296
rect 438308 158244 438360 158296
rect 128176 158176 128228 158228
rect 274364 158176 274416 158228
rect 285404 158176 285456 158228
rect 330576 158176 330628 158228
rect 394240 158176 394292 158228
rect 440608 158176 440660 158228
rect 128728 158108 128780 158160
rect 274456 158108 274508 158160
rect 292304 158108 292356 158160
rect 326436 158108 326488 158160
rect 395896 158108 395948 158160
rect 441896 158108 441948 158160
rect 131488 158040 131540 158092
rect 271696 158040 271748 158092
rect 132408 157972 132460 158024
rect 271604 157972 271656 158024
rect 158536 157904 158588 157956
rect 276020 157904 276072 157956
rect 159916 157836 159968 157888
rect 271328 157836 271380 157888
rect 271420 157836 271472 157888
rect 277952 157836 278004 157888
rect 234620 157768 234672 157820
rect 285496 158040 285548 158092
rect 318156 158040 318208 158092
rect 398472 158040 398524 158092
rect 441804 158040 441856 158092
rect 289360 157972 289412 158024
rect 289544 157972 289596 158024
rect 321652 157972 321704 158024
rect 401048 157972 401100 158024
rect 441712 157972 441764 158024
rect 286140 157904 286192 157956
rect 319444 157904 319496 157956
rect 403992 157904 404044 157956
rect 438216 157904 438268 157956
rect 288256 157836 288308 157888
rect 320548 157836 320600 157888
rect 406476 157836 406528 157888
rect 439688 157836 439740 157888
rect 97632 157632 97684 157684
rect 297364 157632 297416 157684
rect 121920 157564 121972 157616
rect 289360 157564 289412 157616
rect 271328 157496 271380 157548
rect 274640 157496 274692 157548
rect 329748 157428 329800 157480
rect 355232 157428 355284 157480
rect 321560 157360 321612 157412
rect 356980 157360 357032 157412
rect 123208 157292 123260 157344
rect 290740 157292 290792 157344
rect 295708 157292 295760 157344
rect 296352 157292 296404 157344
rect 343916 157292 343968 157344
rect 273720 157224 273772 157276
rect 274180 157224 274232 157276
rect 348700 157224 348752 157276
rect 117320 157156 117372 157208
rect 282736 157156 282788 157208
rect 286876 157156 286928 157208
rect 333612 157156 333664 157208
rect 116492 157088 116544 157140
rect 282828 157088 282880 157140
rect 316040 157088 316092 157140
rect 134892 157020 134944 157072
rect 279976 157020 280028 157072
rect 334532 157020 334584 157072
rect 135904 156952 135956 157004
rect 277216 156952 277268 157004
rect 335636 156952 335688 157004
rect 138112 156884 138164 156936
rect 277124 156884 277176 156936
rect 338120 156884 338172 156936
rect 137008 156816 137060 156868
rect 274548 156816 274600 156868
rect 336832 156816 336884 156868
rect 148876 156748 148928 156800
rect 273720 156748 273772 156800
rect 282736 156748 282788 156800
rect 316960 156748 317012 156800
rect 118240 156680 118292 156732
rect 234620 156680 234672 156732
rect 287428 156680 287480 156732
rect 306380 156680 306432 156732
rect 178868 156612 178920 156664
rect 275376 156612 275428 156664
rect 291936 156612 291988 156664
rect 313280 156612 313332 156664
rect 181812 156544 181864 156596
rect 275284 156544 275336 156596
rect 290740 156544 290792 156596
rect 323124 156544 323176 156596
rect 184020 156476 184072 156528
rect 272524 156476 272576 156528
rect 185952 156408 186004 156460
rect 272616 156408 272668 156460
rect 144092 156340 144144 156392
rect 295708 156340 295760 156392
rect 280068 155864 280120 155916
rect 338212 155864 338264 155916
rect 140688 155796 140740 155848
rect 284116 155796 284168 155848
rect 339500 155796 339552 155848
rect 274640 155728 274692 155780
rect 275836 155728 275888 155780
rect 346676 155728 346728 155780
rect 294328 155660 294380 155712
rect 294972 155660 295024 155712
rect 342352 155660 342404 155712
rect 140504 155592 140556 155644
rect 280068 155592 280120 155644
rect 281448 155592 281500 155644
rect 345112 155592 345164 155644
rect 141792 155524 141844 155576
rect 278596 155524 278648 155576
rect 341064 155524 341116 155576
rect 145288 155456 145340 155508
rect 281448 155456 281500 155508
rect 295708 155456 295760 155508
rect 296536 155456 296588 155508
rect 324228 155456 324280 155508
rect 146392 155388 146444 155440
rect 277308 155388 277360 155440
rect 346400 155388 346452 155440
rect 136088 155320 136140 155372
rect 265716 155320 265768 155372
rect 299296 155320 299348 155372
rect 321560 155320 321612 155372
rect 147680 155252 147732 155304
rect 274640 155252 274692 155304
rect 195888 155184 195940 155236
rect 267004 155184 267056 155236
rect 198464 155116 198516 155168
rect 267188 155116 267240 155168
rect 201040 155048 201092 155100
rect 264336 155048 264388 155100
rect 203432 154980 203484 155032
rect 261576 154980 261628 155032
rect 124588 154912 124640 154964
rect 295708 154912 295760 154964
rect 143080 154844 143132 154896
rect 294328 154844 294380 154896
rect 157064 154776 157116 154828
rect 298376 154776 298428 154828
rect 299296 154776 299348 154828
rect 284760 154572 284812 154624
rect 287428 154572 287480 154624
rect 125416 154504 125468 154556
rect 271788 154504 271840 154556
rect 272708 154504 272760 154556
rect 273168 154504 273220 154556
rect 354404 154504 354456 154556
rect 154120 154436 154172 154488
rect 298008 154436 298060 154488
rect 353300 154436 353352 154488
rect 155776 154368 155828 154420
rect 298560 154368 298612 154420
rect 329748 154368 329800 154420
rect 152648 154300 152700 154352
rect 284208 154300 284260 154352
rect 352196 154300 352248 154352
rect 149888 154232 149940 154284
rect 279884 154232 279936 154284
rect 349804 154232 349856 154284
rect 151360 154164 151412 154216
rect 278688 154164 278740 154216
rect 351000 154164 351052 154216
rect 271788 154096 271840 154148
rect 325332 154096 325384 154148
rect 227720 154028 227772 154080
rect 275008 154028 275060 154080
rect 208400 153960 208452 154012
rect 272340 153960 272392 154012
rect 193220 153892 193272 153944
rect 269672 153892 269724 153944
rect 286048 153892 286100 153944
rect 292948 153892 293000 153944
rect 168380 153824 168432 153876
rect 265440 153824 265492 153876
rect 287336 153824 287388 153876
rect 305000 153824 305052 153876
rect 154488 153756 154540 153808
rect 272708 153756 272760 153808
rect 141424 153144 141476 153196
rect 258908 153144 258960 153196
rect 144368 153076 144420 153128
rect 258816 153076 258868 153128
rect 146024 153008 146076 153060
rect 258724 153008 258776 153060
rect 148508 152940 148560 152992
rect 256148 152940 256200 152992
rect 150992 152872 151044 152924
rect 256240 152872 256292 152924
rect 288900 152668 288952 152720
rect 310520 152668 310572 152720
rect 291660 152600 291712 152652
rect 331220 152600 331272 152652
rect 295616 152532 295668 152584
rect 357440 152532 357492 152584
rect 135260 152464 135312 152516
rect 261484 152464 261536 152516
rect 271236 152464 271288 152516
rect 280436 152464 280488 152516
rect 298192 152464 298244 152516
rect 374092 152464 374144 152516
rect 182180 151104 182232 151156
rect 268200 151104 268252 151156
rect 285956 151104 286008 151156
rect 299572 151104 299624 151156
rect 146300 151036 146352 151088
rect 262588 151036 262640 151088
rect 291568 151036 291620 151088
rect 333980 151036 334032 151088
rect 184940 149812 184992 149864
rect 268108 149812 268160 149864
rect 157340 149744 157392 149796
rect 264152 149744 264204 149796
rect 288808 149744 288860 149796
rect 314660 149744 314712 149796
rect 121460 149676 121512 149728
rect 258448 149676 258500 149728
rect 292856 149676 292908 149728
rect 340880 149676 340932 149728
rect 224960 148384 225012 148436
rect 273904 148384 273956 148436
rect 128360 148316 128412 148368
rect 259920 148316 259972 148368
rect 273996 148316 274048 148368
rect 282000 148316 282052 148368
rect 285864 148316 285916 148368
rect 300860 148316 300912 148368
rect 200120 146956 200172 147008
rect 270868 146956 270920 147008
rect 282000 146956 282052 147008
rect 283380 146956 283432 147008
rect 139400 146888 139452 146940
rect 261392 146888 261444 146940
rect 270960 146888 271012 146940
rect 281908 146888 281960 146940
rect 287244 146888 287296 146940
rect 303620 146888 303672 146940
rect 218060 145664 218112 145716
rect 273536 145664 273588 145716
rect 150440 145596 150492 145648
rect 262496 145596 262548 145648
rect 133880 145528 133932 145580
rect 261300 145528 261352 145580
rect 273904 145528 273956 145580
rect 280344 145528 280396 145580
rect 288716 145528 288768 145580
rect 317420 145528 317472 145580
rect 216680 144304 216732 144356
rect 273444 144304 273496 144356
rect 186320 144236 186372 144288
rect 269580 144236 269632 144288
rect 132500 144168 132552 144220
rect 259828 144168 259880 144220
rect 260196 144168 260248 144220
rect 279148 144168 279200 144220
rect 291476 144168 291528 144220
rect 328460 144168 328512 144220
rect 209780 142944 209832 142996
rect 272248 142944 272300 142996
rect 197360 142876 197412 142928
rect 270776 142876 270828 142928
rect 286324 142876 286376 142928
rect 291476 142876 291528 142928
rect 143540 142808 143592 142860
rect 260104 142808 260156 142860
rect 291384 142808 291436 142860
rect 332600 142808 332652 142860
rect 201500 141516 201552 141568
rect 270684 141516 270736 141568
rect 126980 141448 127032 141500
rect 259736 141448 259788 141500
rect 115940 141380 115992 141432
rect 258356 141380 258408 141432
rect 291292 141380 291344 141432
rect 335360 141380 335412 141432
rect 211160 140156 211212 140208
rect 272156 140156 272208 140208
rect 161480 140088 161532 140140
rect 265348 140088 265400 140140
rect 107660 140020 107712 140072
rect 257068 140020 257120 140072
rect 292764 140020 292816 140072
rect 339500 140020 339552 140072
rect 165620 138728 165672 138780
rect 265256 138728 265308 138780
rect 110420 138660 110472 138712
rect 256976 138660 257028 138712
rect 274088 138660 274140 138712
rect 281816 138660 281868 138712
rect 292672 138660 292724 138712
rect 342260 138660 342312 138712
rect 3516 137912 3568 137964
rect 84844 137912 84896 137964
rect 226340 137300 226392 137352
rect 274916 137300 274968 137352
rect 103520 137232 103572 137284
rect 255688 137232 255740 137284
rect 155960 135872 156012 135924
rect 264060 135872 264112 135924
rect 179420 134580 179472 134632
rect 268016 134580 268068 134632
rect 143632 134512 143684 134564
rect 262404 134512 262456 134564
rect 267004 134512 267056 134564
rect 280712 134512 280764 134564
rect 287152 134512 287204 134564
rect 307760 134512 307812 134564
rect 183560 133220 183612 133272
rect 267924 133220 267976 133272
rect 151820 133152 151872 133204
rect 263968 133152 264020 133204
rect 268568 133152 268620 133204
rect 279056 133152 279108 133204
rect 288624 133152 288676 133204
rect 318800 133152 318852 133204
rect 187700 131792 187752 131844
rect 265624 131792 265676 131844
rect 190460 131724 190512 131776
rect 269488 131724 269540 131776
rect 293316 131724 293368 131776
rect 332692 131724 332744 131776
rect 205640 130500 205692 130552
rect 272064 130500 272116 130552
rect 193312 130432 193364 130484
rect 269396 130432 269448 130484
rect 120080 130364 120132 130416
rect 258264 130364 258316 130416
rect 292580 130364 292632 130416
rect 340972 130364 341024 130416
rect 198740 129072 198792 129124
rect 270592 129072 270644 129124
rect 129740 129004 129792 129056
rect 259644 129004 259696 129056
rect 296168 129004 296220 129056
rect 350540 129004 350592 129056
rect 204260 127644 204312 127696
rect 271144 127644 271196 127696
rect 118700 127576 118752 127628
rect 254584 127576 254636 127628
rect 218152 126284 218204 126336
rect 273352 126284 273404 126336
rect 180800 126216 180852 126268
rect 267832 126216 267884 126268
rect 229100 124924 229152 124976
rect 274824 124924 274876 124976
rect 169760 124856 169812 124908
rect 266728 124856 266780 124908
rect 275284 124856 275336 124908
rect 281724 124856 281776 124908
rect 136640 123428 136692 123480
rect 261208 123428 261260 123480
rect 140780 122068 140832 122120
rect 261116 122068 261168 122120
rect 147680 120708 147732 120760
rect 262312 120708 262364 120760
rect 154580 119348 154632 119400
rect 263876 119348 263928 119400
rect 158720 117920 158772 117972
rect 263784 117920 263836 117972
rect 127072 116560 127124 116612
rect 259552 116560 259604 116612
rect 162860 115200 162912 115252
rect 265164 115200 265216 115252
rect 167000 113772 167052 113824
rect 265072 113772 265124 113824
rect 442264 113092 442316 113144
rect 579804 113092 579856 113144
rect 173900 112412 173952 112464
rect 266636 112412 266688 112464
rect 3148 111732 3200 111784
rect 86224 111732 86276 111784
rect 185032 111052 185084 111104
rect 267740 111052 267792 111104
rect 269856 111052 269908 111104
rect 280528 111052 280580 111104
rect 191840 109692 191892 109744
rect 269304 109692 269356 109744
rect 131120 108264 131172 108316
rect 259460 108264 259512 108316
rect 260104 108264 260156 108316
rect 278964 108264 279016 108316
rect 201592 106904 201644 106956
rect 270500 106904 270552 106956
rect 219440 105612 219492 105664
rect 273260 105612 273312 105664
rect 124220 105544 124272 105596
rect 258172 105544 258224 105596
rect 230480 104184 230532 104236
rect 274732 104184 274784 104236
rect 106280 104116 106332 104168
rect 255596 104116 255648 104168
rect 135352 102756 135404 102808
rect 261024 102756 261076 102808
rect 138020 101396 138072 101448
rect 260932 101396 260984 101448
rect 149060 99968 149112 100020
rect 262772 99968 262824 100020
rect 151912 98608 151964 98660
rect 263692 98608 263744 98660
rect 3516 97928 3568 97980
rect 10324 97928 10376 97980
rect 114560 95888 114612 95940
rect 256884 95888 256936 95940
rect 4804 94460 4856 94512
rect 238760 94460 238812 94512
rect 102140 93100 102192 93152
rect 255504 93100 255556 93152
rect 111800 91740 111852 91792
rect 256792 91740 256844 91792
rect 122840 90312 122892 90364
rect 258540 90312 258592 90364
rect 241612 89224 241664 89276
rect 277860 89224 277912 89276
rect 238760 89156 238812 89208
rect 276204 89156 276256 89208
rect 236000 89088 236052 89140
rect 276296 89088 276348 89140
rect 233240 89020 233292 89072
rect 276388 89020 276440 89072
rect 290280 89020 290332 89072
rect 322940 89020 322992 89072
rect 99380 88952 99432 89004
rect 247776 88952 247828 89004
rect 255504 88952 255556 89004
rect 278044 88952 278096 89004
rect 290188 88952 290240 89004
rect 325700 88952 325752 89004
rect 278964 88748 279016 88800
rect 283288 88748 283340 88800
rect 45560 87592 45612 87644
rect 246396 87592 246448 87644
rect 117320 86232 117372 86284
rect 238024 86232 238076 86284
rect 3516 85484 3568 85536
rect 95884 85484 95936 85536
rect 287060 51688 287112 51740
rect 307852 51688 307904 51740
rect 494704 33056 494756 33108
rect 580172 33056 580224 33108
rect 24860 28228 24912 28280
rect 243268 28228 243320 28280
rect 113180 26868 113232 26920
rect 257160 26868 257212 26920
rect 110512 25508 110564 25560
rect 242164 25508 242216 25560
rect 102232 24080 102284 24132
rect 247684 24080 247736 24132
rect 88340 22720 88392 22772
rect 246304 22720 246356 22772
rect 247408 22720 247460 22772
rect 277768 22720 277820 22772
rect 290096 22720 290148 22772
rect 324320 22720 324372 22772
rect 160100 21360 160152 21412
rect 264520 21360 264572 21412
rect 142160 19932 142212 19984
rect 260840 19932 260892 19984
rect 212540 18572 212592 18624
rect 271972 18572 272024 18624
rect 291200 18572 291252 18624
rect 329840 18572 329892 18624
rect 267740 17280 267792 17332
rect 281632 17280 281684 17332
rect 194600 17212 194652 17264
rect 269212 17212 269264 17264
rect 259460 15852 259512 15904
rect 279516 15852 279568 15904
rect 119896 14424 119948 14476
rect 253204 14424 253256 14476
rect 256700 14424 256752 14476
rect 278872 14424 278924 14476
rect 288532 14424 288584 14476
rect 312176 14424 312228 14476
rect 109040 13064 109092 13116
rect 255964 13064 256016 13116
rect 184940 11772 184992 11824
rect 186136 11772 186188 11824
rect 105728 11704 105780 11756
rect 255412 11704 255464 11756
rect 278044 11568 278096 11620
rect 283196 11568 283248 11620
rect 227536 10344 227588 10396
rect 275100 10344 275152 10396
rect 274824 10276 274876 10328
rect 280804 10276 280856 10328
rect 298100 10276 298152 10328
rect 376024 10276 376076 10328
rect 294604 9188 294656 9240
rect 344560 9188 344612 9240
rect 294236 9120 294288 9172
rect 348056 9120 348108 9172
rect 296076 9052 296128 9104
rect 355232 9052 355284 9104
rect 299388 8984 299440 9036
rect 397736 8984 397788 9036
rect 87972 8916 88024 8968
rect 252928 8916 252980 8968
rect 284668 8916 284720 8968
rect 292488 8916 292540 8968
rect 295064 8916 295116 8968
rect 414296 8916 414348 8968
rect 177856 7624 177908 7676
rect 266544 7624 266596 7676
rect 295524 7624 295576 7676
rect 39580 7556 39632 7608
rect 246028 7556 246080 7608
rect 299572 7556 299624 7608
rect 300768 7556 300820 7608
rect 361120 7556 361172 7608
rect 261760 6876 261812 6928
rect 269764 6876 269816 6928
rect 284576 6876 284628 6928
rect 288992 6876 289044 6928
rect 3424 6808 3476 6860
rect 14464 6808 14516 6860
rect 288440 6808 288492 6860
rect 316224 6808 316276 6860
rect 290004 6740 290056 6792
rect 322112 6740 322164 6792
rect 242900 6672 242952 6724
rect 277676 6672 277728 6724
rect 294144 6672 294196 6724
rect 350448 6672 350500 6724
rect 234620 6604 234672 6656
rect 276572 6604 276624 6656
rect 294052 6604 294104 6656
rect 354036 6604 354088 6656
rect 235816 6536 235868 6588
rect 276112 6536 276164 6588
rect 295432 6536 295484 6588
rect 357532 6536 357584 6588
rect 176660 6468 176712 6520
rect 257344 6468 257396 6520
rect 285772 6468 285824 6520
rect 294880 6468 294932 6520
rect 296720 6468 296772 6520
rect 365812 6468 365864 6520
rect 173164 6400 173216 6452
rect 266452 6400 266504 6452
rect 290648 6400 290700 6452
rect 400128 6400 400180 6452
rect 101036 6332 101088 6384
rect 255780 6332 255832 6384
rect 286968 6332 287020 6384
rect 403624 6332 403676 6384
rect 70308 6264 70360 6316
rect 250260 6264 250312 6316
rect 293592 6264 293644 6316
rect 410800 6264 410852 6316
rect 52552 6196 52604 6248
rect 247316 6196 247368 6248
rect 254676 6196 254728 6248
rect 279240 6196 279292 6248
rect 289728 6196 289780 6248
rect 408408 6196 408460 6248
rect 45468 6128 45520 6180
rect 244924 6128 244976 6180
rect 248788 6128 248840 6180
rect 277584 6128 277636 6180
rect 288348 6128 288400 6180
rect 407212 6128 407264 6180
rect 293316 5448 293368 5500
rect 297272 5448 297324 5500
rect 210976 5244 211028 5296
rect 268384 5244 268436 5296
rect 207388 5176 207440 5228
rect 272432 5176 272484 5228
rect 297364 5176 297416 5228
rect 189724 5108 189776 5160
rect 269948 5108 270000 5160
rect 289820 5108 289872 5160
rect 169576 5040 169628 5092
rect 266912 5040 266964 5092
rect 285680 5040 285732 5092
rect 298468 5040 298520 5092
rect 164884 4972 164936 5024
rect 265532 4972 265584 5024
rect 289912 4972 289964 5024
rect 297364 4972 297416 5024
rect 97448 4904 97500 4956
rect 254124 4904 254176 4956
rect 265348 4904 265400 4956
rect 279424 4904 279476 4956
rect 324412 4972 324464 5024
rect 328000 5040 328052 5092
rect 48964 4836 49016 4888
rect 247224 4836 247276 4888
rect 15936 4768 15988 4820
rect 241980 4768 242032 4820
rect 245200 4768 245252 4820
rect 277492 4836 277544 4888
rect 293960 4836 294012 4888
rect 349252 4836 349304 4888
rect 295340 4768 295392 4820
rect 359924 4768 359976 4820
rect 278688 4360 278740 4412
rect 282092 4360 282144 4412
rect 287704 4156 287756 4208
rect 290188 4156 290240 4208
rect 12348 4088 12400 4140
rect 18604 4088 18656 4140
rect 253480 4088 253532 4140
rect 260196 4088 260248 4140
rect 285588 4088 285640 4140
rect 338672 4088 338724 4140
rect 429660 4088 429712 4140
rect 440516 4088 440568 4140
rect 292396 4020 292448 4072
rect 297456 4020 297508 4072
rect 298744 4020 298796 4072
rect 369400 4020 369452 4072
rect 427268 4020 427320 4072
rect 437848 4020 437900 4072
rect 6460 3952 6512 4004
rect 7656 3952 7708 4004
rect 295248 3952 295300 4004
rect 384764 3952 384816 4004
rect 426164 3952 426216 4004
rect 437480 3952 437532 4004
rect 266544 3884 266596 3936
rect 269856 3884 269908 3936
rect 293868 3884 293920 3936
rect 391848 3884 391900 3936
rect 423772 3884 423824 3936
rect 437664 3884 437716 3936
rect 5264 3816 5316 3868
rect 7564 3816 7616 3868
rect 171968 3816 172020 3868
rect 239404 3816 239456 3868
rect 293776 3816 293828 3868
rect 395344 3816 395396 3868
rect 424968 3816 425020 3868
rect 439136 3816 439188 3868
rect 460204 3816 460256 3868
rect 462780 3816 462832 3868
rect 516784 3816 516836 3868
rect 519544 3816 519596 3868
rect 566464 3816 566516 3868
rect 569132 3816 569184 3868
rect 135260 3748 135312 3800
rect 136456 3748 136508 3800
rect 161296 3748 161348 3800
rect 264244 3748 264296 3800
rect 294972 3748 295024 3800
rect 125876 3680 125928 3732
rect 238116 3680 238168 3732
rect 244096 3680 244148 3732
rect 278136 3680 278188 3732
rect 296628 3680 296680 3732
rect 298100 3748 298152 3800
rect 398932 3748 398984 3800
rect 422576 3748 422628 3800
rect 438952 3748 439004 3800
rect 2872 3544 2924 3596
rect 13084 3612 13136 3664
rect 28908 3612 28960 3664
rect 39304 3612 39356 3664
rect 43076 3612 43128 3664
rect 57244 3612 57296 3664
rect 7656 3544 7708 3596
rect 572 3476 624 3528
rect 4804 3476 4856 3528
rect 9956 3476 10008 3528
rect 11704 3476 11756 3528
rect 20628 3544 20680 3596
rect 68284 3612 68336 3664
rect 93952 3612 94004 3664
rect 254400 3612 254452 3664
rect 264152 3612 264204 3664
rect 273904 3612 273956 3664
rect 291108 3612 291160 3664
rect 402520 3680 402572 3732
rect 421380 3680 421432 3732
rect 438032 3680 438084 3732
rect 67916 3544 67968 3596
rect 71044 3544 71096 3596
rect 77300 3544 77352 3596
rect 78220 3544 78272 3596
rect 85672 3544 85724 3596
rect 88984 3544 89036 3596
rect 90364 3544 90416 3596
rect 254308 3544 254360 3596
rect 262956 3544 263008 3596
rect 267004 3544 267056 3596
rect 267096 3544 267148 3596
rect 271236 3544 271288 3596
rect 283012 3544 283064 3596
rect 284300 3544 284352 3596
rect 285036 3544 285088 3596
rect 17224 3476 17276 3528
rect 21824 3476 21876 3528
rect 22744 3476 22796 3528
rect 24216 3476 24268 3528
rect 4068 3408 4120 3460
rect 4896 3408 4948 3460
rect 11152 3408 11204 3460
rect 30104 3476 30156 3528
rect 31024 3476 31076 3528
rect 33600 3476 33652 3528
rect 35164 3476 35216 3528
rect 38384 3476 38436 3528
rect 39396 3476 39448 3528
rect 51356 3476 51408 3528
rect 247684 3476 247736 3528
rect 251180 3476 251232 3528
rect 268568 3476 268620 3528
rect 268844 3476 268896 3528
rect 274088 3476 274140 3528
rect 277124 3476 277176 3528
rect 282184 3476 282236 3528
rect 32404 3408 32456 3460
rect 35992 3408 36044 3460
rect 50344 3408 50396 3460
rect 43444 3340 43496 3392
rect 47860 3340 47912 3392
rect 247132 3408 247184 3460
rect 249984 3408 250036 3460
rect 268476 3408 268528 3460
rect 270040 3408 270092 3460
rect 273996 3408 274048 3460
rect 276020 3408 276072 3460
rect 291844 3476 291896 3528
rect 296076 3476 296128 3528
rect 409604 3612 409656 3664
rect 420184 3612 420236 3664
rect 438860 3612 438912 3664
rect 297456 3544 297508 3596
rect 406016 3544 406068 3596
rect 418988 3544 419040 3596
rect 437572 3544 437624 3596
rect 442356 3544 442408 3596
rect 447416 3544 447468 3596
rect 453304 3544 453356 3596
rect 455696 3544 455748 3596
rect 467104 3544 467156 3596
rect 469864 3544 469916 3596
rect 475384 3544 475436 3596
rect 476948 3544 477000 3596
rect 500224 3544 500276 3596
rect 501788 3544 501840 3596
rect 511264 3544 511316 3596
rect 513564 3544 513616 3596
rect 413100 3476 413152 3528
rect 417884 3476 417936 3528
rect 439228 3476 439280 3528
rect 440332 3476 440384 3528
rect 441528 3476 441580 3528
rect 448612 3476 448664 3528
rect 449808 3476 449860 3528
rect 462964 3476 463016 3528
rect 465172 3476 465224 3528
rect 538864 3476 538916 3528
rect 540796 3476 540848 3528
rect 547880 3476 547932 3528
rect 548708 3476 548760 3528
rect 556160 3476 556212 3528
rect 556988 3476 557040 3528
rect 563704 3476 563756 3528
rect 565636 3476 565688 3528
rect 571984 3476 572036 3528
rect 573916 3476 573968 3528
rect 581000 3476 581052 3528
rect 581828 3476 581880 3528
rect 292304 3408 292356 3460
rect 416688 3408 416740 3460
rect 60740 3340 60792 3392
rect 61660 3340 61712 3392
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 260656 3340 260708 3392
rect 267096 3340 267148 3392
rect 295984 3340 296036 3392
rect 346952 3340 347004 3392
rect 357440 3340 357492 3392
rect 358728 3340 358780 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 415492 3340 415544 3392
rect 439044 3408 439096 3460
rect 445116 3408 445168 3460
rect 458088 3408 458140 3460
rect 458824 3408 458876 3460
rect 484032 3408 484084 3460
rect 514116 3408 514168 3460
rect 514760 3408 514812 3460
rect 527916 3408 527968 3460
rect 533712 3408 533764 3460
rect 570604 3408 570656 3460
rect 572720 3408 572772 3460
rect 428464 3340 428516 3392
rect 437756 3340 437808 3392
rect 446404 3340 446456 3392
rect 452108 3340 452160 3392
rect 514024 3340 514076 3392
rect 515956 3340 516008 3392
rect 554044 3340 554096 3392
rect 559748 3340 559800 3392
rect 17040 3272 17092 3324
rect 21364 3272 21416 3324
rect 293500 3272 293552 3324
rect 298100 3272 298152 3324
rect 307760 3272 307812 3324
rect 309048 3272 309100 3324
rect 324320 3272 324372 3324
rect 325608 3272 325660 3324
rect 332692 3272 332744 3324
rect 333888 3272 333940 3324
rect 340880 3272 340932 3324
rect 342168 3272 342220 3324
rect 430856 3272 430908 3324
rect 439320 3272 439372 3324
rect 504364 3272 504416 3324
rect 507676 3272 507728 3324
rect 1676 3204 1728 3256
rect 8944 3204 8996 3256
rect 252376 3204 252428 3256
rect 260104 3204 260156 3256
rect 272432 3204 272484 3256
rect 275284 3204 275336 3256
rect 432052 3204 432104 3256
rect 439504 3204 439556 3256
rect 280712 3136 280764 3188
rect 283196 3136 283248 3188
rect 476764 3136 476816 3188
rect 479340 3136 479392 3188
rect 485044 3136 485096 3188
rect 487620 3136 487672 3188
rect 534724 3136 534776 3188
rect 537208 3136 537260 3188
rect 560944 3136 560996 3188
rect 563244 3136 563296 3188
rect 567844 3136 567896 3188
rect 570328 3136 570380 3188
rect 471244 3068 471296 3120
rect 473452 3068 473504 3120
rect 520924 3068 520976 3120
rect 523040 3068 523092 3120
rect 284484 3000 284536 3052
rect 286600 3000 286652 3052
rect 464344 3000 464396 3052
rect 466276 3000 466328 3052
rect 478236 3000 478288 3052
rect 480536 3000 480588 3052
rect 503076 3000 503128 3052
rect 505376 3000 505428 3052
rect 8760 2932 8812 2984
rect 10416 2932 10468 2984
rect 19432 2932 19484 2984
rect 25504 2932 25556 2984
rect 457444 2932 457496 2984
rect 459192 2932 459244 2984
rect 494796 2864 494848 2916
rect 499396 2864 499448 2916
rect 273628 2796 273680 2848
rect 278688 2796 278740 2848
rect 316040 1096 316092 1148
rect 317328 1096 317380 1148
<< obsm1 >>
rect 220000 480000 356620 563308
rect 100000 160000 236620 243308
rect 300000 160000 436620 243308
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 2832 632088 2834 632097
rect 2778 632023 2834 632032
rect 3330 606112 3386 606121
rect 3330 606047 3386 606056
rect 3344 605878 3372 606047
rect 3332 605872 3384 605878
rect 3332 605814 3384 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3146 553888 3202 553897
rect 3146 553823 3202 553832
rect 3160 553722 3188 553823
rect 3148 553716 3200 553722
rect 3148 553658 3200 553664
rect 3330 527912 3386 527921
rect 3330 527847 3386 527856
rect 3344 527202 3372 527847
rect 3332 527196 3384 527202
rect 3332 527138 3384 527144
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 2870 501800 2926 501809
rect 2870 501735 2926 501744
rect 2884 501022 2912 501735
rect 2872 501016 2924 501022
rect 2872 500958 2924 500964
rect 3330 475688 3386 475697
rect 3330 475623 3386 475632
rect 3344 474774 3372 475623
rect 3332 474768 3384 474774
rect 3332 474710 3384 474716
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3344 462398 3372 462567
rect 3332 462392 3384 462398
rect 3332 462334 3384 462340
rect 2870 449576 2926 449585
rect 2870 449511 2926 449520
rect 2884 447846 2912 449511
rect 3436 449342 3464 671191
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 4804 632120 4856 632126
rect 4804 632062 4856 632068
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3424 449336 3476 449342
rect 3424 449278 3476 449284
rect 3528 449274 3556 619103
rect 3606 566944 3662 566953
rect 3606 566879 3662 566888
rect 3516 449268 3568 449274
rect 3516 449210 3568 449216
rect 3620 449206 3648 566879
rect 4816 465730 4844 632062
rect 6932 474026 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 21364 656940 21416 656946
rect 21364 656882 21416 656888
rect 17224 605872 17276 605878
rect 17224 605814 17276 605820
rect 10324 579692 10376 579698
rect 10324 579634 10376 579640
rect 8944 553716 8996 553722
rect 8944 553658 8996 553664
rect 6920 474020 6972 474026
rect 6920 473962 6972 473968
rect 4804 465724 4856 465730
rect 4804 465666 4856 465672
rect 8956 460222 8984 553658
rect 10336 469878 10364 579634
rect 14464 527196 14516 527202
rect 14464 527138 14516 527144
rect 13084 501016 13136 501022
rect 13084 500958 13136 500964
rect 10324 469872 10376 469878
rect 10324 469814 10376 469820
rect 8944 460216 8996 460222
rect 8944 460158 8996 460164
rect 13096 457502 13124 500958
rect 14476 471306 14504 527138
rect 17236 472666 17264 605814
rect 18604 514820 18656 514826
rect 18604 514762 18656 514768
rect 17224 472660 17276 472666
rect 17224 472602 17276 472608
rect 14464 471300 14516 471306
rect 14464 471242 14516 471248
rect 13084 457496 13136 457502
rect 13084 457438 13136 457444
rect 18616 456074 18644 514762
rect 21376 478174 21404 656882
rect 21364 478168 21416 478174
rect 21364 478110 21416 478116
rect 18604 456068 18656 456074
rect 18604 456010 18656 456016
rect 23492 449410 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 40052 461650 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40040 461644 40092 461650
rect 40040 461586 40092 461592
rect 23480 449404 23532 449410
rect 23480 449346 23532 449352
rect 3608 449200 3660 449206
rect 3608 449142 3660 449148
rect 71792 447914 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 88352 449478 88380 702406
rect 105464 699786 105492 703520
rect 105452 699780 105504 699786
rect 105452 699722 105504 699728
rect 108304 699780 108356 699786
rect 108304 699722 108356 699728
rect 108316 468518 108344 699722
rect 108304 468512 108356 468518
rect 108304 468454 108356 468460
rect 88340 449472 88392 449478
rect 88340 449414 88392 449420
rect 136652 447982 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 153212 449614 153240 702406
rect 169772 464370 169800 702406
rect 171784 683188 171836 683194
rect 171784 683130 171836 683136
rect 171796 467158 171824 683130
rect 171784 467152 171836 467158
rect 171784 467094 171836 467100
rect 169760 464364 169812 464370
rect 169760 464306 169812 464312
rect 153200 449608 153252 449614
rect 153200 449550 153252 449556
rect 201512 448118 201540 702986
rect 217968 700324 218020 700330
rect 217968 700266 218020 700272
rect 217874 516896 217930 516905
rect 217874 516831 217930 516840
rect 217782 515944 217838 515953
rect 217782 515879 217838 515888
rect 217690 513768 217746 513777
rect 217690 513703 217746 513712
rect 217598 489968 217654 489977
rect 217598 489903 217654 489912
rect 217506 488336 217562 488345
rect 217506 488271 217562 488280
rect 217322 488064 217378 488073
rect 217322 487999 217378 488008
rect 217336 478922 217364 487999
rect 217324 478916 217376 478922
rect 217324 478858 217376 478864
rect 217520 476814 217548 488271
rect 217508 476808 217560 476814
rect 217508 476750 217560 476756
rect 217612 451926 217640 489903
rect 217704 472734 217732 513703
rect 217692 472728 217744 472734
rect 217692 472670 217744 472676
rect 217796 471374 217824 515879
rect 217784 471368 217836 471374
rect 217784 471310 217836 471316
rect 217888 454714 217916 516831
rect 217876 454708 217928 454714
rect 217876 454650 217928 454656
rect 217600 451920 217652 451926
rect 217600 451862 217652 451868
rect 201500 448112 201552 448118
rect 201500 448054 201552 448060
rect 136640 447976 136692 447982
rect 136640 447918 136692 447924
rect 71780 447908 71832 447914
rect 71780 447850 71832 447856
rect 2872 447840 2924 447846
rect 2872 447782 2924 447788
rect 217980 446758 218008 700266
rect 218072 478242 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 235184 700330 235212 703520
rect 267660 700330 267688 703520
rect 283852 700398 283880 703520
rect 300136 700466 300164 703520
rect 332520 700534 332548 703520
rect 348804 700602 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700596 348844 700602
rect 348792 700538 348844 700544
rect 357716 700596 357768 700602
rect 357716 700538 357768 700544
rect 332508 700528 332560 700534
rect 332508 700470 332560 700476
rect 300124 700460 300176 700466
rect 300124 700402 300176 700408
rect 357624 700460 357676 700466
rect 357624 700402 357676 700408
rect 283840 700392 283892 700398
rect 283840 700334 283892 700340
rect 357532 700392 357584 700398
rect 357532 700334 357584 700340
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 357440 700324 357492 700330
rect 357440 700266 357492 700272
rect 219346 512816 219402 512825
rect 219346 512751 219402 512760
rect 219162 511048 219218 511057
rect 219162 510983 219218 510992
rect 219070 508192 219126 508201
rect 219070 508127 219126 508136
rect 218060 478236 218112 478242
rect 218060 478178 218112 478184
rect 219084 475386 219112 508127
rect 219072 475380 219124 475386
rect 219072 475322 219124 475328
rect 219176 474094 219204 510983
rect 219254 509960 219310 509969
rect 219254 509895 219310 509904
rect 219164 474088 219216 474094
rect 219164 474030 219216 474036
rect 219268 458862 219296 509895
rect 219256 458856 219308 458862
rect 219256 458798 219308 458804
rect 219360 450566 219388 512751
rect 220084 478916 220136 478922
rect 220084 478858 220136 478864
rect 219348 450560 219400 450566
rect 219348 450502 219400 450508
rect 217968 446752 218020 446758
rect 217968 446694 218020 446700
rect 220096 446486 220124 478858
rect 309140 478304 309192 478310
rect 309140 478246 309192 478252
rect 242898 477320 242954 477329
rect 242898 477255 242954 477264
rect 233332 476808 233384 476814
rect 233332 476750 233384 476756
rect 220084 446480 220136 446486
rect 220084 446422 220136 446428
rect 230940 446004 230992 446010
rect 230940 445946 230992 445952
rect 229744 445936 229796 445942
rect 229744 445878 229796 445884
rect 10324 445800 10376 445806
rect 10324 445742 10376 445748
rect 7564 444440 7616 444446
rect 7564 444382 7616 444388
rect 3516 443692 3568 443698
rect 3516 443634 3568 443640
rect 3424 442264 3476 442270
rect 3424 442206 3476 442212
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 3332 411256 3384 411262
rect 3332 411198 3384 411204
rect 3344 410553 3372 411198
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3332 398812 3384 398818
rect 3332 398754 3384 398760
rect 3344 397497 3372 398754
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3056 372564 3108 372570
rect 3056 372506 3108 372512
rect 3068 371385 3096 372506
rect 3054 371376 3110 371385
rect 3054 371311 3110 371320
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3332 320136 3384 320142
rect 3332 320078 3384 320084
rect 3344 319297 3372 320078
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3332 293956 3384 293962
rect 3332 293898 3384 293904
rect 3344 293185 3372 293898
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 2964 267708 3016 267714
rect 2964 267650 3016 267656
rect 2976 267209 3004 267650
rect 2962 267200 3018 267209
rect 2962 267135 3018 267144
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3240 241460 3292 241466
rect 3240 241402 3292 241408
rect 3252 241097 3280 241402
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3148 189032 3200 189038
rect 3148 188974 3200 188980
rect 3160 188873 3188 188974
rect 3146 188864 3202 188873
rect 3146 188799 3202 188808
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3436 45529 3464 442206
rect 3528 201929 3556 443634
rect 3608 440904 3660 440910
rect 3608 440846 3660 440852
rect 3620 358465 3648 440846
rect 7576 423638 7604 444382
rect 7564 423632 7616 423638
rect 7564 423574 7616 423580
rect 3606 358456 3662 358465
rect 3606 358391 3662 358400
rect 7564 308440 7616 308446
rect 7564 308382 7616 308388
rect 4896 280832 4948 280838
rect 4896 280774 4948 280780
rect 3608 244928 3660 244934
rect 3608 244870 3660 244876
rect 3514 201920 3570 201929
rect 3514 201855 3570 201864
rect 3516 164212 3568 164218
rect 3516 164154 3568 164160
rect 3528 162897 3556 164154
rect 3514 162888 3570 162897
rect 3514 162823 3570 162832
rect 3620 149841 3648 244870
rect 3606 149832 3662 149841
rect 3606 149767 3662 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 4804 94512 4856 94518
rect 4804 94454 4856 94460
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 584 480 612 3470
rect 1676 3256 1728 3262
rect 1676 3198 1728 3204
rect 1688 480 1716 3198
rect 2884 480 2912 3538
rect 4816 3534 4844 94454
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4908 3466 4936 280774
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 5264 3868 5316 3874
rect 5264 3810 5316 3816
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4080 480 4108 3402
rect 5276 480 5304 3810
rect 6472 480 6500 3946
rect 7576 3874 7604 308382
rect 8944 307080 8996 307086
rect 8944 307022 8996 307028
rect 7656 265668 7708 265674
rect 7656 265610 7708 265616
rect 7668 4010 7696 265610
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7564 3868 7616 3874
rect 7564 3810 7616 3816
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7668 480 7696 3538
rect 8956 3262 8984 307022
rect 10336 97986 10364 445742
rect 228456 445188 228508 445194
rect 228456 445130 228508 445136
rect 225604 444984 225656 444990
rect 225604 444926 225656 444932
rect 224224 444848 224276 444854
rect 224224 444790 224276 444796
rect 95976 444712 96028 444718
rect 95976 444654 96028 444660
rect 93124 444644 93176 444650
rect 93124 444586 93176 444592
rect 86224 444576 86276 444582
rect 86224 444518 86276 444524
rect 84844 444508 84896 444514
rect 84844 444450 84896 444456
rect 14464 443012 14516 443018
rect 14464 442954 14516 442960
rect 13084 304292 13136 304298
rect 13084 304234 13136 304240
rect 12440 294636 12492 294642
rect 12440 294578 12492 294584
rect 10416 279472 10468 279478
rect 10416 279414 10468 279420
rect 10324 97980 10376 97986
rect 10324 97922 10376 97928
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 8944 3256 8996 3262
rect 8944 3198 8996 3204
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8772 480 8800 2926
rect 9968 480 9996 3470
rect 10428 2990 10456 279414
rect 11704 260160 11756 260166
rect 11704 260102 11756 260108
rect 11716 3534 11744 260102
rect 12452 16574 12480 294578
rect 12452 16546 13032 16574
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 11164 480 11192 3402
rect 12360 480 12388 4082
rect 13004 3482 13032 16546
rect 13096 3670 13124 304234
rect 13820 250504 13872 250510
rect 13820 250446 13872 250452
rect 13832 16574 13860 250446
rect 13832 16546 14320 16574
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 13004 3454 13584 3482
rect 13556 480 13584 3454
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 14476 6866 14504 442954
rect 39304 309120 39356 309126
rect 39304 309062 39356 309068
rect 32404 308644 32456 308650
rect 32404 308586 32456 308592
rect 25504 308508 25556 308514
rect 25504 308450 25556 308456
rect 18604 304360 18656 304366
rect 18604 304302 18656 304308
rect 17224 302932 17276 302938
rect 17224 302874 17276 302880
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 15948 480 15976 4762
rect 17236 3534 17264 302874
rect 17960 264240 18012 264246
rect 17960 264182 18012 264188
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17040 3324 17092 3330
rect 17040 3266 17092 3272
rect 17052 480 17080 3266
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 264182
rect 18616 4146 18644 304302
rect 21364 300144 21416 300150
rect 21364 300086 21416 300092
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19444 480 19472 2926
rect 20640 480 20668 3538
rect 21376 3330 21404 300086
rect 22744 298784 22796 298790
rect 22744 298726 22796 298732
rect 22100 290488 22152 290494
rect 22100 290430 22152 290436
rect 22112 16574 22140 290430
rect 22112 16546 22600 16574
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 21364 3324 21416 3330
rect 21364 3266 21416 3272
rect 21836 480 21864 3470
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 22756 3534 22784 298726
rect 24860 28280 24912 28286
rect 24860 28222 24912 28228
rect 24872 16574 24900 28222
rect 24872 16546 25360 16574
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24228 480 24256 3470
rect 25332 480 25360 16546
rect 25516 2990 25544 308450
rect 31024 307148 31076 307154
rect 31024 307090 31076 307096
rect 27620 303000 27672 303006
rect 27620 302942 27672 302948
rect 26240 284980 26292 284986
rect 26240 284922 26292 284928
rect 25504 2984 25556 2990
rect 25504 2926 25556 2932
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 284922
rect 27632 16574 27660 302942
rect 30380 289128 30432 289134
rect 30380 289070 30432 289076
rect 30392 16574 30420 289070
rect 27632 16546 27752 16574
rect 30392 16546 30880 16574
rect 27724 480 27752 16546
rect 28908 3664 28960 3670
rect 28908 3606 28960 3612
rect 28920 480 28948 3606
rect 30104 3528 30156 3534
rect 30104 3470 30156 3476
rect 30116 480 30144 3470
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31036 3534 31064 307090
rect 31760 247716 31812 247722
rect 31760 247658 31812 247664
rect 31772 16574 31800 247658
rect 31772 16546 31984 16574
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 32416 3466 32444 308586
rect 35164 305652 35216 305658
rect 35164 305594 35216 305600
rect 34520 287700 34572 287706
rect 34520 287642 34572 287648
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 33612 480 33640 3470
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 287642
rect 35176 3534 35204 305594
rect 35900 297424 35952 297430
rect 35900 297366 35952 297372
rect 35912 16574 35940 297366
rect 35912 16546 36768 16574
rect 35164 3528 35216 3534
rect 35164 3470 35216 3476
rect 35992 3460 36044 3466
rect 35992 3402 36044 3408
rect 36004 480 36032 3402
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 39316 3670 39344 309062
rect 68284 308916 68336 308922
rect 68284 308858 68336 308864
rect 57244 308848 57296 308854
rect 57244 308790 57296 308796
rect 50344 308780 50396 308786
rect 50344 308722 50396 308728
rect 43444 308712 43496 308718
rect 43444 308654 43496 308660
rect 39396 301504 39448 301510
rect 39396 301446 39448 301452
rect 39304 3664 39356 3670
rect 39304 3606 39356 3612
rect 39408 3534 39436 301446
rect 40040 283620 40092 283626
rect 40040 283562 40092 283568
rect 40052 16574 40080 283562
rect 41420 262880 41472 262886
rect 41420 262822 41472 262828
rect 41432 16574 41460 262822
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 39580 7608 39632 7614
rect 39580 7550 39632 7556
rect 38384 3528 38436 3534
rect 38384 3470 38436 3476
rect 39396 3528 39448 3534
rect 39396 3470 39448 3476
rect 38396 480 38424 3470
rect 39592 480 39620 7550
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 43076 3664 43128 3670
rect 43076 3606 43128 3612
rect 43088 480 43116 3606
rect 43456 3398 43484 308654
rect 49700 286340 49752 286346
rect 49700 286282 49752 286288
rect 44180 282192 44232 282198
rect 44180 282134 44232 282140
rect 44192 16574 44220 282134
rect 45560 87644 45612 87650
rect 45560 87586 45612 87592
rect 45572 16574 45600 87586
rect 49712 16574 49740 286282
rect 44192 16546 44312 16574
rect 45572 16546 46704 16574
rect 49712 16546 50200 16574
rect 43444 3392 43496 3398
rect 43444 3334 43496 3340
rect 44284 480 44312 16546
rect 45468 6180 45520 6186
rect 45468 6122 45520 6128
rect 45480 480 45508 6122
rect 46676 480 46704 16546
rect 48964 4888 49016 4894
rect 48964 4830 49016 4836
rect 47860 3392 47912 3398
rect 47860 3334 47912 3340
rect 47872 480 47900 3334
rect 48976 480 49004 4830
rect 50172 480 50200 16546
rect 50356 3466 50384 308722
rect 52460 307216 52512 307222
rect 52460 307158 52512 307164
rect 52472 16574 52500 307158
rect 53840 298852 53892 298858
rect 53840 298794 53892 298800
rect 53852 16574 53880 298794
rect 55220 275324 55272 275330
rect 55220 275266 55272 275272
rect 55232 16574 55260 275266
rect 56600 258732 56652 258738
rect 56600 258674 56652 258680
rect 56612 16574 56640 258674
rect 52472 16546 53328 16574
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 52552 6248 52604 6254
rect 52552 6190 52604 6196
rect 51356 3528 51408 3534
rect 51356 3470 51408 3476
rect 50344 3460 50396 3466
rect 50344 3402 50396 3408
rect 51368 480 51396 3470
rect 52564 480 52592 6190
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 57256 3670 57284 308790
rect 64880 307284 64932 307290
rect 64880 307226 64932 307232
rect 57980 297492 58032 297498
rect 57980 297434 58032 297440
rect 57992 16574 58020 297434
rect 60740 295996 60792 296002
rect 60740 295938 60792 295944
rect 59360 273964 59412 273970
rect 59360 273906 59412 273912
rect 57992 16546 58480 16574
rect 57244 3664 57296 3670
rect 57244 3606 57296 3612
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 273906
rect 60752 3398 60780 295938
rect 63500 285048 63552 285054
rect 63500 284990 63552 284996
rect 62120 272536 62172 272542
rect 62120 272478 62172 272484
rect 60832 253224 60884 253230
rect 60832 253166 60884 253172
rect 60740 3392 60792 3398
rect 60740 3334 60792 3340
rect 60844 480 60872 253166
rect 62132 16574 62160 272478
rect 63512 16574 63540 284990
rect 64892 16574 64920 307226
rect 66260 271176 66312 271182
rect 66260 271118 66312 271124
rect 66272 16574 66300 271118
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 64892 16546 65104 16574
rect 66272 16546 66760 16574
rect 61660 3392 61712 3398
rect 61660 3334 61712 3340
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61672 354 61700 3334
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66732 480 66760 16546
rect 68296 3670 68324 308858
rect 71780 305720 71832 305726
rect 71780 305662 71832 305668
rect 71044 300212 71096 300218
rect 71044 300154 71096 300160
rect 70400 298920 70452 298926
rect 70400 298862 70452 298868
rect 69020 294704 69072 294710
rect 69020 294646 69072 294652
rect 69032 16574 69060 294646
rect 70412 16574 70440 298862
rect 69032 16546 69152 16574
rect 70412 16546 70992 16574
rect 68284 3664 68336 3670
rect 68284 3606 68336 3612
rect 67916 3596 67968 3602
rect 67916 3538 67968 3544
rect 67928 480 67956 3538
rect 69124 480 69152 16546
rect 70308 6316 70360 6322
rect 70308 6258 70360 6264
rect 70320 480 70348 6258
rect 70964 3482 70992 16546
rect 71056 3602 71084 300154
rect 71792 16574 71820 305662
rect 82820 303068 82872 303074
rect 82820 303010 82872 303016
rect 80060 296064 80112 296070
rect 80060 296006 80112 296012
rect 75920 291848 75972 291854
rect 75920 291790 75972 291796
rect 73160 269816 73212 269822
rect 73160 269758 73212 269764
rect 73172 16574 73200 269758
rect 74540 251864 74592 251870
rect 74540 251806 74592 251812
rect 74552 16574 74580 251806
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 71044 3596 71096 3602
rect 71044 3538 71096 3544
rect 70964 3454 71544 3482
rect 71516 480 71544 3454
rect 72620 480 72648 16546
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 291790
rect 78680 290556 78732 290562
rect 78680 290498 78732 290504
rect 77300 283688 77352 283694
rect 77300 283630 77352 283636
rect 77312 3602 77340 283630
rect 77392 268388 77444 268394
rect 77392 268330 77444 268336
rect 77300 3596 77352 3602
rect 77300 3538 77352 3544
rect 77404 480 77432 268330
rect 78692 16574 78720 290498
rect 80072 16574 80100 296006
rect 81440 282260 81492 282266
rect 81440 282202 81492 282208
rect 81452 16574 81480 282202
rect 82832 16574 82860 303010
rect 84200 265736 84252 265742
rect 84200 265678 84252 265684
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 78220 3596 78272 3602
rect 78220 3538 78272 3544
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78232 354 78260 3538
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 265678
rect 84856 137970 84884 444450
rect 85580 289196 85632 289202
rect 85580 289138 85632 289144
rect 84844 137964 84896 137970
rect 84844 137906 84896 137912
rect 85592 16574 85620 289138
rect 86236 111790 86264 444518
rect 88984 305788 89036 305794
rect 88984 305730 89036 305736
rect 86224 111784 86276 111790
rect 86224 111726 86276 111732
rect 88340 22772 88392 22778
rect 88340 22714 88392 22720
rect 88352 16574 88380 22714
rect 85592 16546 86448 16574
rect 88352 16546 88932 16574
rect 85672 3596 85724 3602
rect 85672 3538 85724 3544
rect 85684 480 85712 3538
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 87972 8968 88024 8974
rect 87972 8910 88024 8916
rect 87984 480 88012 8910
rect 88904 3482 88932 16546
rect 88996 3602 89024 305730
rect 91100 304428 91152 304434
rect 91100 304370 91152 304376
rect 91112 16574 91140 304370
rect 92480 297560 92532 297566
rect 92480 297502 92532 297508
rect 91112 16546 91600 16574
rect 88984 3596 89036 3602
rect 88984 3538 89036 3544
rect 90364 3596 90416 3602
rect 90364 3538 90416 3544
rect 88904 3454 89208 3482
rect 89180 480 89208 3454
rect 90376 480 90404 3538
rect 91572 480 91600 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 86838 -960 86950 326
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92492 354 92520 297502
rect 93136 164218 93164 444586
rect 95884 443148 95936 443154
rect 95884 443090 95936 443096
rect 94504 443080 94556 443086
rect 94504 443022 94556 443028
rect 93860 293276 93912 293282
rect 93860 293218 93912 293224
rect 93124 164212 93176 164218
rect 93124 164154 93176 164160
rect 93872 16574 93900 293218
rect 94516 189038 94544 443022
rect 95240 246356 95292 246362
rect 95240 246298 95292 246304
rect 94504 189032 94556 189038
rect 94504 188974 94556 188980
rect 95252 16574 95280 246298
rect 95896 85542 95924 443090
rect 95988 215286 96016 444654
rect 157984 443284 158036 443290
rect 157984 443226 158036 443232
rect 97264 443216 97316 443222
rect 97264 443158 97316 443164
rect 97276 241466 97304 443158
rect 97906 305688 97962 305697
rect 97906 305623 97962 305632
rect 97724 243500 97776 243506
rect 97724 243442 97776 243448
rect 97264 241460 97316 241466
rect 97264 241402 97316 241408
rect 95976 215280 96028 215286
rect 95976 215222 96028 215228
rect 97736 196897 97764 243442
rect 97816 243432 97868 243438
rect 97816 243374 97868 243380
rect 97722 196888 97778 196897
rect 97722 196823 97778 196832
rect 97828 195945 97856 243374
rect 97814 195936 97870 195945
rect 97814 195871 97870 195880
rect 97814 193760 97870 193769
rect 97814 193695 97870 193704
rect 97722 192808 97778 192817
rect 97722 192743 97778 192752
rect 97538 191040 97594 191049
rect 97538 190975 97594 190984
rect 97446 188184 97502 188193
rect 97446 188119 97502 188128
rect 97354 169960 97410 169969
rect 97354 169895 97410 169904
rect 97368 159594 97396 169895
rect 97460 159934 97488 188119
rect 97448 159928 97500 159934
rect 97448 159870 97500 159876
rect 97552 159866 97580 190975
rect 97630 189952 97686 189961
rect 97630 189887 97686 189896
rect 97540 159860 97592 159866
rect 97540 159802 97592 159808
rect 97356 159588 97408 159594
rect 97356 159530 97408 159536
rect 97644 157690 97672 189887
rect 97736 159798 97764 192743
rect 97724 159792 97776 159798
rect 97724 159734 97776 159740
rect 97828 159730 97856 193695
rect 97920 168473 97948 305623
rect 98000 291916 98052 291922
rect 98000 291858 98052 291864
rect 97906 168464 97962 168473
rect 97906 168399 97962 168408
rect 97906 168328 97962 168337
rect 97906 168263 97962 168272
rect 97816 159724 97868 159730
rect 97816 159666 97868 159672
rect 97920 159662 97948 168263
rect 97908 159656 97960 159662
rect 97908 159598 97960 159604
rect 97632 157684 97684 157690
rect 97632 157626 97684 157632
rect 95884 85536 95936 85542
rect 95884 85478 95936 85484
rect 98012 16574 98040 291858
rect 157996 255270 158024 443226
rect 224236 293962 224264 444790
rect 224224 293956 224276 293962
rect 224224 293898 224276 293904
rect 225616 267714 225644 444926
rect 228364 443488 228416 443494
rect 228364 443430 228416 443436
rect 228376 306338 228404 443430
rect 228468 320142 228496 445130
rect 228548 443556 228600 443562
rect 228548 443498 228600 443504
rect 228560 411262 228588 443498
rect 228548 411256 228600 411262
rect 228548 411198 228600 411204
rect 228456 320136 228508 320142
rect 228456 320078 228508 320084
rect 228364 306332 228416 306338
rect 228364 306274 228416 306280
rect 225604 267708 225656 267714
rect 225604 267650 225656 267656
rect 157984 255264 158036 255270
rect 157984 255206 158036 255212
rect 229756 244934 229784 445878
rect 230846 445768 230902 445777
rect 230846 445703 230902 445712
rect 229928 445120 229980 445126
rect 229928 445062 229980 445068
rect 229836 443420 229888 443426
rect 229836 443362 229888 443368
rect 229848 346390 229876 443362
rect 229940 372570 229968 445062
rect 230020 444916 230072 444922
rect 230020 444858 230072 444864
rect 230032 398818 230060 444858
rect 230860 442270 230888 445703
rect 230848 442264 230900 442270
rect 230848 442206 230900 442212
rect 230952 440910 230980 445946
rect 233344 443306 233372 476750
rect 238760 476604 238812 476610
rect 238760 476546 238812 476552
rect 236000 476536 236052 476542
rect 236000 476478 236052 476484
rect 235906 476232 235962 476241
rect 235906 476167 235962 476176
rect 235920 476134 235948 476167
rect 234620 476128 234672 476134
rect 234620 476070 234672 476076
rect 235908 476128 235960 476134
rect 235908 476070 235960 476076
rect 234632 447030 234660 476070
rect 234712 451920 234764 451926
rect 234712 451862 234764 451868
rect 234620 447024 234672 447030
rect 234620 446966 234672 446972
rect 234344 446480 234396 446486
rect 234344 446422 234396 446428
rect 233344 443278 233634 443306
rect 234356 443292 234384 446422
rect 234724 443306 234752 451862
rect 235540 447024 235592 447030
rect 235540 446966 235592 446972
rect 235552 443306 235580 446966
rect 236012 443612 236040 476478
rect 236092 476468 236144 476474
rect 236092 476410 236144 476416
rect 236104 460934 236132 476410
rect 237286 476368 237342 476377
rect 237286 476303 237288 476312
rect 237340 476303 237342 476312
rect 237288 476274 237340 476280
rect 237378 476232 237434 476241
rect 237378 476167 237434 476176
rect 237392 460934 237420 476167
rect 236104 460906 236960 460934
rect 237392 460906 237696 460934
rect 236012 443584 236224 443612
rect 236196 443306 236224 443584
rect 236932 443306 236960 460906
rect 237668 443306 237696 460906
rect 238772 447030 238800 476546
rect 242912 476542 242940 477255
rect 255226 477048 255282 477057
rect 255226 476983 255282 476992
rect 264978 477048 265034 477057
rect 264978 476983 265034 476992
rect 270498 477048 270554 477057
rect 270498 476983 270554 476992
rect 304998 477048 305054 477057
rect 304998 476983 305054 476992
rect 307758 477048 307814 477057
rect 307758 476983 307814 476992
rect 251180 476740 251232 476746
rect 251180 476682 251232 476688
rect 244278 476640 244334 476649
rect 244278 476575 244280 476584
rect 244332 476575 244334 476584
rect 247038 476640 247094 476649
rect 247038 476575 247094 476584
rect 244280 476546 244332 476552
rect 242900 476536 242952 476542
rect 242900 476478 242952 476484
rect 242992 476536 243044 476542
rect 242992 476478 243044 476484
rect 238852 476332 238904 476338
rect 238852 476274 238904 476280
rect 240140 476332 240192 476338
rect 240140 476274 240192 476280
rect 238760 447024 238812 447030
rect 238760 446966 238812 446972
rect 238864 443306 238892 476274
rect 239220 447024 239272 447030
rect 239220 446966 239272 446972
rect 234724 443278 235106 443306
rect 235552 443278 235842 443306
rect 236196 443278 236578 443306
rect 236932 443278 237314 443306
rect 237668 443278 238050 443306
rect 238786 443278 238892 443306
rect 239232 443306 239260 446966
rect 240152 443306 240180 476274
rect 241520 476264 241572 476270
rect 240230 476232 240286 476241
rect 240230 476167 240286 476176
rect 241426 476232 241482 476241
rect 241520 476206 241572 476212
rect 242806 476232 242862 476241
rect 241426 476167 241482 476176
rect 240244 460934 240272 476167
rect 241440 476134 241468 476167
rect 241428 476128 241480 476134
rect 241428 476070 241480 476076
rect 240244 460906 240640 460934
rect 240612 443306 240640 460906
rect 241532 447030 241560 476206
rect 243004 476218 243032 476478
rect 247052 476474 247080 476575
rect 248420 476536 248472 476542
rect 248420 476478 248472 476484
rect 249890 476504 249946 476513
rect 247040 476468 247092 476474
rect 247040 476410 247092 476416
rect 245752 476400 245804 476406
rect 244278 476368 244334 476377
rect 245752 476342 245804 476348
rect 244278 476303 244334 476312
rect 244292 476270 244320 476303
rect 242806 476167 242808 476176
rect 242860 476167 242862 476176
rect 242912 476190 243032 476218
rect 244280 476264 244332 476270
rect 244280 476206 244332 476212
rect 245658 476232 245714 476241
rect 244924 476196 244976 476202
rect 242808 476138 242860 476144
rect 241612 475380 241664 475386
rect 241612 475322 241664 475328
rect 241520 447024 241572 447030
rect 241520 446966 241572 446972
rect 241624 443306 241652 475322
rect 242164 447024 242216 447030
rect 242164 446966 242216 446972
rect 242176 443306 242204 446966
rect 242912 443306 242940 476190
rect 245658 476167 245714 476176
rect 244924 476138 244976 476144
rect 242992 476128 243044 476134
rect 242992 476070 243044 476076
rect 244280 476128 244332 476134
rect 244280 476070 244332 476076
rect 243004 460934 243032 476070
rect 243004 460906 243584 460934
rect 243556 443306 243584 460906
rect 244292 447030 244320 476070
rect 244372 458856 244424 458862
rect 244372 458798 244424 458804
rect 244280 447024 244332 447030
rect 244280 446966 244332 446972
rect 244384 443306 244412 458798
rect 244936 446282 244964 476138
rect 245672 476134 245700 476167
rect 245660 476128 245712 476134
rect 245660 476070 245712 476076
rect 245108 447024 245160 447030
rect 245108 446966 245160 446972
rect 244924 446276 244976 446282
rect 244924 446218 244976 446224
rect 245120 443306 245148 446966
rect 245764 443306 245792 476342
rect 247222 476232 247278 476241
rect 247222 476167 247278 476176
rect 247132 474088 247184 474094
rect 247132 474030 247184 474036
rect 246856 446276 246908 446282
rect 246856 446218 246908 446224
rect 239232 443278 239522 443306
rect 240152 443278 240258 443306
rect 240612 443278 240994 443306
rect 241624 443278 241730 443306
rect 242176 443278 242466 443306
rect 242912 443278 243202 443306
rect 243556 443278 243938 443306
rect 244384 443278 244674 443306
rect 245120 443278 245410 443306
rect 245764 443278 246146 443306
rect 246868 443292 246896 446218
rect 247144 443306 247172 474030
rect 247236 460934 247264 476167
rect 248432 460934 248460 476478
rect 249890 476439 249946 476448
rect 249904 476270 249932 476439
rect 249892 476264 249944 476270
rect 249798 476232 249854 476241
rect 249892 476206 249944 476212
rect 249798 476167 249854 476176
rect 249812 460934 249840 476167
rect 247236 460906 248000 460934
rect 248432 460906 248736 460934
rect 249812 460906 250208 460934
rect 247972 443306 248000 460906
rect 248708 443306 248736 460906
rect 249800 450560 249852 450566
rect 249800 450502 249852 450508
rect 247144 443278 247618 443306
rect 247972 443278 248354 443306
rect 248708 443278 249090 443306
rect 249812 443292 249840 450502
rect 250180 443306 250208 460906
rect 251088 446072 251140 446078
rect 251088 446014 251140 446020
rect 251100 443698 251128 446014
rect 251088 443692 251140 443698
rect 251088 443634 251140 443640
rect 251192 443306 251220 476682
rect 255240 476678 255268 476983
rect 255318 476912 255374 476921
rect 255318 476847 255374 476856
rect 255228 476672 255280 476678
rect 252558 476640 252614 476649
rect 255228 476614 255280 476620
rect 252558 476575 252560 476584
rect 252612 476575 252614 476584
rect 252652 476604 252704 476610
rect 252560 476546 252612 476552
rect 252652 476546 252704 476552
rect 252466 476368 252522 476377
rect 252466 476303 252522 476312
rect 251822 476232 251878 476241
rect 251822 476167 251878 476176
rect 251272 472728 251324 472734
rect 251272 472670 251324 472676
rect 251284 460934 251312 472670
rect 251284 460906 251680 460934
rect 251652 443306 251680 460906
rect 251836 447030 251864 476167
rect 252480 476134 252508 476303
rect 252468 476128 252520 476134
rect 252468 476070 252520 476076
rect 252664 460934 252692 476546
rect 255332 476406 255360 476847
rect 264992 476814 265020 476983
rect 255412 476808 255464 476814
rect 264980 476808 265032 476814
rect 255412 476750 255464 476756
rect 260838 476776 260894 476785
rect 255320 476400 255372 476406
rect 255320 476342 255372 476348
rect 253202 476232 253258 476241
rect 253202 476167 253258 476176
rect 254582 476232 254638 476241
rect 254582 476167 254638 476176
rect 252664 460906 253152 460934
rect 251824 447024 251876 447030
rect 251824 446966 251876 446972
rect 252744 447024 252796 447030
rect 252744 446966 252796 446972
rect 250180 443278 250562 443306
rect 251192 443278 251298 443306
rect 251652 443278 252034 443306
rect 252756 443292 252784 446966
rect 253124 443306 253152 460906
rect 253216 446554 253244 476167
rect 253940 476128 253992 476134
rect 253940 476070 253992 476076
rect 253952 447030 253980 476070
rect 254032 471368 254084 471374
rect 254032 471310 254084 471316
rect 253940 447024 253992 447030
rect 253940 446966 253992 446972
rect 253204 446548 253256 446554
rect 253204 446490 253256 446496
rect 254044 443306 254072 471310
rect 254596 447098 254624 476167
rect 255424 470594 255452 476750
rect 264980 476750 265032 476756
rect 260838 476711 260840 476720
rect 260892 476711 260894 476720
rect 260840 476682 260892 476688
rect 259460 476672 259512 476678
rect 258078 476640 258134 476649
rect 258078 476575 258134 476584
rect 258262 476640 258318 476649
rect 259460 476614 259512 476620
rect 263598 476640 263654 476649
rect 258262 476575 258318 476584
rect 256792 476468 256844 476474
rect 256792 476410 256844 476416
rect 256606 476232 256662 476241
rect 256606 476167 256662 476176
rect 255332 470566 255452 470594
rect 254584 447092 254636 447098
rect 254584 447034 254636 447040
rect 254676 447024 254728 447030
rect 254676 446966 254728 446972
rect 254688 443306 254716 446966
rect 255332 443306 255360 470566
rect 256056 454708 256108 454714
rect 256056 454650 256108 454656
rect 256068 443306 256096 454650
rect 256620 446486 256648 476167
rect 256804 460934 256832 476410
rect 258092 476406 258120 476575
rect 258276 476542 258304 476575
rect 258264 476536 258316 476542
rect 258264 476478 258316 476484
rect 258080 476400 258132 476406
rect 258080 476342 258132 476348
rect 258172 476332 258224 476338
rect 258172 476274 258224 476280
rect 257986 476232 258042 476241
rect 257986 476167 258042 476176
rect 256804 460906 257568 460934
rect 257160 446548 257212 446554
rect 257160 446490 257212 446496
rect 256608 446480 256660 446486
rect 256608 446422 256660 446428
rect 253124 443278 253506 443306
rect 254044 443278 254242 443306
rect 254688 443278 254978 443306
rect 255332 443278 255714 443306
rect 256068 443278 256450 443306
rect 257172 443292 257200 446490
rect 257540 443306 257568 460906
rect 258000 446554 258028 476167
rect 258184 460934 258212 476274
rect 259472 460934 259500 476614
rect 263598 476575 263600 476584
rect 263652 476575 263654 476584
rect 263600 476546 263652 476552
rect 262312 476536 262364 476542
rect 262312 476478 262364 476484
rect 267922 476504 267978 476513
rect 260104 476400 260156 476406
rect 260932 476400 260984 476406
rect 260104 476342 260156 476348
rect 260746 476368 260802 476377
rect 258184 460906 259040 460934
rect 259472 460906 259776 460934
rect 258632 447092 258684 447098
rect 258632 447034 258684 447040
rect 257988 446548 258040 446554
rect 257988 446490 258040 446496
rect 257540 443278 257922 443306
rect 258644 443292 258672 447034
rect 259012 443306 259040 460906
rect 259748 443306 259776 460906
rect 260116 446962 260144 476342
rect 260932 476342 260984 476348
rect 260746 476303 260802 476312
rect 260760 476134 260788 476303
rect 260748 476128 260800 476134
rect 260748 476070 260800 476076
rect 260104 446956 260156 446962
rect 260104 446898 260156 446904
rect 260944 443306 260972 476342
rect 261482 476232 261538 476241
rect 261482 476167 261538 476176
rect 262126 476232 262182 476241
rect 262126 476167 262128 476176
rect 261496 447030 261524 476167
rect 262180 476167 262182 476176
rect 262128 476138 262180 476144
rect 261484 447024 261536 447030
rect 261484 446966 261536 446972
rect 261576 446480 261628 446486
rect 261576 446422 261628 446428
rect 259012 443278 259394 443306
rect 259748 443278 260130 443306
rect 260866 443278 260972 443306
rect 261588 443292 261616 446422
rect 262324 443292 262352 476478
rect 267922 476439 267924 476448
rect 267976 476439 267978 476448
rect 267924 476410 267976 476416
rect 267646 476368 267702 476377
rect 267646 476303 267702 476312
rect 263692 476264 263744 476270
rect 263506 476232 263562 476241
rect 263692 476206 263744 476212
rect 264886 476232 264942 476241
rect 263506 476167 263562 476176
rect 263520 476134 263548 476167
rect 262864 476128 262916 476134
rect 262864 476070 262916 476076
rect 263508 476128 263560 476134
rect 263508 476070 263560 476076
rect 262876 447098 262904 476070
rect 262864 447092 262916 447098
rect 262864 447034 262916 447040
rect 263048 446548 263100 446554
rect 263048 446490 263100 446496
rect 263060 443292 263088 446490
rect 263704 443306 263732 476206
rect 264244 476196 264296 476202
rect 264886 476167 264942 476176
rect 266266 476232 266322 476241
rect 266266 476167 266322 476176
rect 267554 476232 267610 476241
rect 267554 476167 267610 476176
rect 264244 476138 264296 476144
rect 264256 446894 264284 476138
rect 264900 451926 264928 476167
rect 265624 476128 265676 476134
rect 265624 476070 265676 476076
rect 265072 456136 265124 456142
rect 265072 456078 265124 456084
rect 264888 451920 264940 451926
rect 264888 451862 264940 451868
rect 264520 446956 264572 446962
rect 264520 446898 264572 446904
rect 264244 446888 264296 446894
rect 264244 446830 264296 446836
rect 263704 443278 263810 443306
rect 264532 443292 264560 446898
rect 265084 443306 265112 456078
rect 265636 446962 265664 476070
rect 266280 450566 266308 476167
rect 266452 457564 266504 457570
rect 266452 457506 266504 457512
rect 266268 450560 266320 450566
rect 266268 450502 266320 450508
rect 265992 447024 266044 447030
rect 265992 446966 266044 446972
rect 265624 446956 265676 446962
rect 265624 446898 265676 446904
rect 265084 443278 265282 443306
rect 266004 443292 266032 446966
rect 266464 443306 266492 457506
rect 267568 454714 267596 476167
rect 267556 454708 267608 454714
rect 267556 454650 267608 454656
rect 267660 453354 267688 476303
rect 270512 476270 270540 476983
rect 277858 476912 277914 476921
rect 277858 476847 277914 476856
rect 277584 476740 277636 476746
rect 277584 476682 277636 476688
rect 276018 476640 276074 476649
rect 276018 476575 276074 476584
rect 276032 476542 276060 476575
rect 276020 476536 276072 476542
rect 273258 476504 273314 476513
rect 276020 476478 276072 476484
rect 273258 476439 273314 476448
rect 273272 476406 273300 476439
rect 273260 476400 273312 476406
rect 273260 476342 273312 476348
rect 274454 476368 274510 476377
rect 274454 476303 274510 476312
rect 270500 476264 270552 476270
rect 269026 476232 269082 476241
rect 269026 476167 269082 476176
rect 270406 476232 270462 476241
rect 270500 476206 270552 476212
rect 271786 476232 271842 476241
rect 270406 476167 270462 476176
rect 271786 476167 271842 476176
rect 273166 476232 273222 476241
rect 273166 476167 273222 476176
rect 267832 469940 267884 469946
rect 267832 469882 267884 469888
rect 267648 453348 267700 453354
rect 267648 453290 267700 453296
rect 267464 447092 267516 447098
rect 267464 447034 267516 447040
rect 266464 443278 266754 443306
rect 267476 443292 267504 447034
rect 267844 443306 267872 469882
rect 269040 452062 269068 476167
rect 269212 468580 269264 468586
rect 269212 468522 269264 468528
rect 269224 460934 269252 468522
rect 269224 460906 269344 460934
rect 269028 452056 269080 452062
rect 269028 451998 269080 452004
rect 268936 446956 268988 446962
rect 268936 446898 268988 446904
rect 267844 443278 268226 443306
rect 268948 443292 268976 446898
rect 269316 443306 269344 460906
rect 270420 450702 270448 476167
rect 270776 460284 270828 460290
rect 270776 460226 270828 460232
rect 270408 450696 270460 450702
rect 270408 450638 270460 450644
rect 270408 447092 270460 447098
rect 270408 447034 270460 447040
rect 269316 443278 269698 443306
rect 270420 443292 270448 447034
rect 270788 443306 270816 460226
rect 271800 453490 271828 476167
rect 273180 458930 273208 476167
rect 273168 458924 273220 458930
rect 273168 458866 273220 458872
rect 274468 454850 274496 476303
rect 274546 476232 274602 476241
rect 274546 476167 274602 476176
rect 275926 476232 275982 476241
rect 275926 476167 275982 476176
rect 277306 476232 277362 476241
rect 277306 476167 277362 476176
rect 274456 454844 274508 454850
rect 274456 454786 274508 454792
rect 271788 453484 271840 453490
rect 271788 453426 271840 453432
rect 271880 451920 271932 451926
rect 271880 451862 271932 451868
rect 272248 451920 272300 451926
rect 272248 451862 272300 451868
rect 270788 443278 271170 443306
rect 271892 443292 271920 451862
rect 272260 443306 272288 451862
rect 274088 450628 274140 450634
rect 274088 450570 274140 450576
rect 273352 450560 273404 450566
rect 273352 450502 273404 450508
rect 272260 443278 272642 443306
rect 273364 443292 273392 450502
rect 274100 443292 274128 450570
rect 274560 450566 274588 476167
rect 274640 453348 274692 453354
rect 274640 453290 274692 453296
rect 275192 453348 275244 453354
rect 275192 453290 275244 453296
rect 274548 450560 274600 450566
rect 274548 450502 274600 450508
rect 274652 443306 274680 453290
rect 275204 443306 275232 453290
rect 275940 451994 275968 476167
rect 276020 454776 276072 454782
rect 276020 454718 276072 454724
rect 275928 451988 275980 451994
rect 275928 451930 275980 451936
rect 276032 447030 276060 454718
rect 276112 454708 276164 454714
rect 276112 454650 276164 454656
rect 276020 447024 276072 447030
rect 276020 446966 276072 446972
rect 276124 443306 276152 454650
rect 277320 453422 277348 476167
rect 277596 460934 277624 476682
rect 277872 476134 277900 476847
rect 302238 476776 302294 476785
rect 302238 476711 302240 476720
rect 302292 476711 302294 476720
rect 302240 476682 302292 476688
rect 305012 476678 305040 476983
rect 278780 476672 278832 476678
rect 278780 476614 278832 476620
rect 305000 476672 305052 476678
rect 305000 476614 305052 476620
rect 278686 476232 278742 476241
rect 278686 476167 278742 476176
rect 277860 476128 277912 476134
rect 277860 476070 277912 476076
rect 277596 460906 278176 460934
rect 277308 453416 277360 453422
rect 277308 453358 277360 453364
rect 277492 452056 277544 452062
rect 277492 451998 277544 452004
rect 276756 447024 276808 447030
rect 276756 446966 276808 446972
rect 276768 443306 276796 446966
rect 277504 443306 277532 451998
rect 278148 443306 278176 460906
rect 278700 458862 278728 476167
rect 278792 460934 278820 476614
rect 282920 476604 282972 476610
rect 282920 476546 282972 476552
rect 280160 476536 280212 476542
rect 280160 476478 280212 476484
rect 280066 476232 280122 476241
rect 280066 476167 280122 476176
rect 278792 460906 279648 460934
rect 278688 458856 278740 458862
rect 278688 458798 278740 458804
rect 279240 450696 279292 450702
rect 279240 450638 279292 450644
rect 274652 443278 274850 443306
rect 275204 443278 275586 443306
rect 276124 443278 276322 443306
rect 276768 443278 277058 443306
rect 277504 443278 277794 443306
rect 278148 443278 278530 443306
rect 279252 443292 279280 450638
rect 279620 443306 279648 460906
rect 280080 454714 280108 476167
rect 280068 454708 280120 454714
rect 280068 454650 280120 454656
rect 280172 447030 280200 476478
rect 280250 476232 280306 476241
rect 280250 476167 280306 476176
rect 280264 456142 280292 476167
rect 281816 458924 281868 458930
rect 281816 458866 281868 458872
rect 280252 456136 280304 456142
rect 280252 456078 280304 456084
rect 280344 453484 280396 453490
rect 280344 453426 280396 453432
rect 280160 447024 280212 447030
rect 280160 446966 280212 446972
rect 280356 443306 280384 453426
rect 281172 447024 281224 447030
rect 281172 446966 281224 446972
rect 281184 443306 281212 446966
rect 281828 443306 281856 458866
rect 279620 443278 280002 443306
rect 280356 443278 280738 443306
rect 281184 443278 281474 443306
rect 281828 443278 282210 443306
rect 282932 443292 282960 476546
rect 307772 476542 307800 476983
rect 307760 476536 307812 476542
rect 307760 476478 307812 476484
rect 285680 476468 285732 476474
rect 285680 476410 285732 476416
rect 284300 476400 284352 476406
rect 284300 476342 284352 476348
rect 283010 476232 283066 476241
rect 283010 476167 283066 476176
rect 283024 457570 283052 476167
rect 283012 457564 283064 457570
rect 283012 457506 283064 457512
rect 283288 454844 283340 454850
rect 283288 454786 283340 454792
rect 283300 443306 283328 454786
rect 284312 443306 284340 476342
rect 285128 450560 285180 450566
rect 285128 450502 285180 450508
rect 283300 443278 283682 443306
rect 284312 443278 284418 443306
rect 285140 443292 285168 450502
rect 285692 443306 285720 476410
rect 287060 476332 287112 476338
rect 287060 476274 287112 476280
rect 285770 476232 285826 476241
rect 285770 476167 285826 476176
rect 285784 469946 285812 476167
rect 285772 469940 285824 469946
rect 285772 469882 285824 469888
rect 286232 451988 286284 451994
rect 286232 451930 286284 451936
rect 286244 443306 286272 451930
rect 287072 443306 287100 476274
rect 288440 476264 288492 476270
rect 287150 476232 287206 476241
rect 288440 476206 288492 476212
rect 289910 476232 289966 476241
rect 287150 476167 287206 476176
rect 287164 468586 287192 476167
rect 287152 468580 287204 468586
rect 287152 468522 287204 468528
rect 287704 453416 287756 453422
rect 287704 453358 287756 453364
rect 287716 443306 287744 453358
rect 288452 443306 288480 476206
rect 289820 476196 289872 476202
rect 289910 476167 289966 476176
rect 292578 476232 292634 476241
rect 292578 476167 292634 476176
rect 295430 476232 295486 476241
rect 295430 476167 295486 476176
rect 298190 476232 298246 476241
rect 298190 476167 298246 476176
rect 300858 476232 300914 476241
rect 300858 476167 300914 476176
rect 289820 476138 289872 476144
rect 289176 458856 289228 458862
rect 289176 458798 289228 458804
rect 289188 443306 289216 458798
rect 289832 443306 289860 476138
rect 289924 460290 289952 476167
rect 291200 476128 291252 476134
rect 291200 476070 291252 476076
rect 291212 460934 291240 476070
rect 291212 460906 291424 460934
rect 289912 460284 289964 460290
rect 289912 460226 289964 460232
rect 290648 454708 290700 454714
rect 290648 454650 290700 454656
rect 290660 443306 290688 454650
rect 291396 443306 291424 460906
rect 292592 451926 292620 476167
rect 295340 467220 295392 467226
rect 295340 467162 295392 467168
rect 292580 451920 292632 451926
rect 292580 451862 292632 451868
rect 294696 450560 294748 450566
rect 294696 450502 294748 450508
rect 293224 446208 293276 446214
rect 293224 446150 293276 446156
rect 292488 446140 292540 446146
rect 292488 446082 292540 446088
rect 285692 443278 285890 443306
rect 286244 443278 286626 443306
rect 287072 443278 287362 443306
rect 287716 443278 288098 443306
rect 288452 443278 288834 443306
rect 289188 443278 289570 443306
rect 289832 443278 290306 443306
rect 290660 443278 291042 443306
rect 291396 443278 291778 443306
rect 292500 443292 292528 446082
rect 293236 443292 293264 446150
rect 293960 445868 294012 445874
rect 293960 445810 294012 445816
rect 293972 443292 294000 445810
rect 294708 443292 294736 450502
rect 295352 446978 295380 467162
rect 295444 450634 295472 476167
rect 298100 469940 298152 469946
rect 298100 469882 298152 469888
rect 296720 451920 296772 451926
rect 296720 451862 296772 451868
rect 295432 450628 295484 450634
rect 295432 450570 295484 450576
rect 295352 446950 295840 446978
rect 295432 444780 295484 444786
rect 295432 444722 295484 444728
rect 295444 443292 295472 444722
rect 295812 443306 295840 446950
rect 296732 443306 296760 451862
rect 297638 444408 297694 444417
rect 297638 444343 297694 444352
rect 295812 443278 296194 443306
rect 296732 443278 296930 443306
rect 297652 443292 297680 444343
rect 298112 443306 298140 469882
rect 298204 453354 298232 476167
rect 299480 471368 299532 471374
rect 299480 471310 299532 471316
rect 299492 460934 299520 471310
rect 299492 460906 300256 460934
rect 298744 454708 298796 454714
rect 298744 454650 298796 454656
rect 298192 453348 298244 453354
rect 298192 453290 298244 453296
rect 298756 443306 298784 454650
rect 300124 443352 300176 443358
rect 298112 443278 298402 443306
rect 298756 443278 299138 443306
rect 299874 443300 300124 443306
rect 299874 443294 300176 443300
rect 300228 443306 300256 460906
rect 300872 454782 300900 476167
rect 302240 475380 302292 475386
rect 302240 475322 302292 475328
rect 300860 454776 300912 454782
rect 300860 454718 300912 454724
rect 300952 453348 301004 453354
rect 300952 453290 301004 453296
rect 300964 443306 300992 453290
rect 302056 446616 302108 446622
rect 302056 446558 302108 446564
rect 299874 443278 300164 443294
rect 300228 443278 300610 443306
rect 300964 443278 301346 443306
rect 302068 443292 302096 446558
rect 302252 446026 302280 475322
rect 307760 460284 307812 460290
rect 307760 460226 307812 460232
rect 305368 457564 305420 457570
rect 305368 457506 305420 457512
rect 303160 456136 303212 456142
rect 303160 456078 303212 456084
rect 302252 445998 302464 446026
rect 302436 443306 302464 445998
rect 303172 443306 303200 456078
rect 305000 449540 305052 449546
rect 305000 449482 305052 449488
rect 304264 446276 304316 446282
rect 304264 446218 304316 446224
rect 302436 443278 302818 443306
rect 303172 443278 303554 443306
rect 304276 443292 304304 446218
rect 305012 443292 305040 449482
rect 305380 443306 305408 457506
rect 307208 449676 307260 449682
rect 307208 449618 307260 449624
rect 306472 446344 306524 446350
rect 306472 446286 306524 446292
rect 305380 443278 305762 443306
rect 306484 443292 306512 446286
rect 307220 443292 307248 449618
rect 307772 443306 307800 460226
rect 308680 443624 308732 443630
rect 308680 443566 308732 443572
rect 307772 443278 307970 443306
rect 308692 443292 308720 443566
rect 309152 443306 309180 478246
rect 313372 478236 313424 478242
rect 313372 478178 313424 478184
rect 310518 476912 310574 476921
rect 310518 476847 310574 476856
rect 310532 476610 310560 476847
rect 310520 476604 310572 476610
rect 310520 476546 310572 476552
rect 313278 476504 313334 476513
rect 313278 476439 313334 476448
rect 313292 476406 313320 476439
rect 313280 476400 313332 476406
rect 313280 476342 313332 476348
rect 313384 470594 313412 478178
rect 346492 478168 346544 478174
rect 346492 478110 346544 478116
rect 322938 476912 322994 476921
rect 322938 476847 322994 476856
rect 314658 476504 314714 476513
rect 314658 476439 314660 476448
rect 314712 476439 314714 476448
rect 314660 476410 314712 476416
rect 317418 476368 317474 476377
rect 317418 476303 317420 476312
rect 317472 476303 317474 476312
rect 320178 476368 320234 476377
rect 320178 476303 320234 476312
rect 317420 476274 317472 476280
rect 320192 476270 320220 476303
rect 320180 476264 320232 476270
rect 320180 476206 320232 476212
rect 322952 476202 322980 476847
rect 325790 476232 325846 476241
rect 322940 476196 322992 476202
rect 325790 476167 325846 476176
rect 322940 476138 322992 476144
rect 325804 476134 325832 476167
rect 325792 476128 325844 476134
rect 325792 476070 325844 476076
rect 329840 474768 329892 474774
rect 329840 474710 329892 474716
rect 327080 471300 327132 471306
rect 327080 471242 327132 471248
rect 313292 470566 313412 470594
rect 313292 447134 313320 470566
rect 324320 469872 324372 469878
rect 324320 469814 324372 469820
rect 316040 468512 316092 468518
rect 316040 468454 316092 468460
rect 318800 468512 318852 468518
rect 318800 468454 318852 468460
rect 313372 464364 313424 464370
rect 313372 464306 313424 464312
rect 313384 460934 313412 464306
rect 316052 460934 316080 468454
rect 313384 460906 314240 460934
rect 316052 460906 316448 460934
rect 313292 447106 313504 447134
rect 312360 446752 312412 446758
rect 312360 446694 312412 446700
rect 311624 446548 311676 446554
rect 311624 446490 311676 446496
rect 310152 446480 310204 446486
rect 310152 446422 310204 446428
rect 309152 443278 309442 443306
rect 310164 443292 310192 446422
rect 310888 446412 310940 446418
rect 310888 446354 310940 446360
rect 310900 443292 310928 446354
rect 311636 443292 311664 446490
rect 312372 443292 312400 446694
rect 313096 443692 313148 443698
rect 313096 443634 313148 443640
rect 313108 443292 313136 443634
rect 313476 443306 313504 447106
rect 314212 443306 314240 460906
rect 316040 449608 316092 449614
rect 316040 449550 316092 449556
rect 315304 443760 315356 443766
rect 315304 443702 315356 443708
rect 313476 443278 313858 443306
rect 314212 443278 314594 443306
rect 315316 443292 315344 443702
rect 316052 443292 316080 449550
rect 316420 443306 316448 460906
rect 317420 458856 317472 458862
rect 317420 458798 317472 458804
rect 317432 443306 317460 458798
rect 318248 449472 318300 449478
rect 318248 449414 318300 449420
rect 316420 443278 316802 443306
rect 317432 443278 317538 443306
rect 318260 443292 318288 449414
rect 318812 445058 318840 468454
rect 320180 467152 320232 467158
rect 320180 467094 320232 467100
rect 318892 461644 318944 461650
rect 318892 461586 318944 461592
rect 318800 445052 318852 445058
rect 318800 444994 318852 445000
rect 318904 443306 318932 461586
rect 320192 460934 320220 467094
rect 322940 465724 322992 465730
rect 322940 465666 322992 465672
rect 321560 461644 321612 461650
rect 321560 461586 321612 461592
rect 320192 460906 320864 460934
rect 320456 449404 320508 449410
rect 320456 449346 320508 449352
rect 319444 445052 319496 445058
rect 319444 444994 319496 445000
rect 319456 443306 319484 444994
rect 318904 443278 319010 443306
rect 319456 443278 319746 443306
rect 320468 443292 320496 449346
rect 320836 443306 320864 460906
rect 321572 443306 321600 461586
rect 322664 449336 322716 449342
rect 322664 449278 322716 449284
rect 320836 443278 321218 443306
rect 321572 443278 321954 443306
rect 322676 443292 322704 449278
rect 322952 443306 322980 465666
rect 323032 464364 323084 464370
rect 323032 464306 323084 464312
rect 323044 460934 323072 464306
rect 324332 460934 324360 469814
rect 325700 465724 325752 465730
rect 325700 465666 325752 465672
rect 325712 460934 325740 465666
rect 327092 460934 327120 471242
rect 323044 460906 323808 460934
rect 324332 460906 325280 460934
rect 325712 460906 326016 460934
rect 327092 460906 327488 460934
rect 323780 443306 323808 460906
rect 324872 449268 324924 449274
rect 324872 449210 324924 449216
rect 322952 443278 323426 443306
rect 323780 443278 324162 443306
rect 324884 443292 324912 449210
rect 325252 443306 325280 460906
rect 325988 443306 326016 460906
rect 327080 449200 327132 449206
rect 327080 449142 327132 449148
rect 325252 443278 325634 443306
rect 325988 443278 326370 443306
rect 327092 443292 327120 449142
rect 327460 443306 327488 460906
rect 328920 456068 328972 456074
rect 328920 456010 328972 456016
rect 328552 448044 328604 448050
rect 328552 447986 328604 447992
rect 327460 443278 327842 443306
rect 328564 443292 328592 447986
rect 328932 443306 328960 456010
rect 329852 443306 329880 474710
rect 345112 474020 345164 474026
rect 345112 473962 345164 473968
rect 332600 472728 332652 472734
rect 332600 472670 332652 472676
rect 329932 463004 329984 463010
rect 329932 462946 329984 462952
rect 329944 460934 329972 462946
rect 331312 462392 331364 462398
rect 331312 462334 331364 462340
rect 329944 460906 330432 460934
rect 330404 443306 330432 460906
rect 331324 443306 331352 462334
rect 332232 444440 332284 444446
rect 332232 444382 332284 444388
rect 328932 443278 329314 443306
rect 329852 443278 330050 443306
rect 330404 443278 330786 443306
rect 331324 443278 331522 443306
rect 332244 443292 332272 444382
rect 332612 443306 332640 472670
rect 345124 460934 345152 473962
rect 346504 460934 346532 478110
rect 347780 472660 347832 472666
rect 347780 472602 347832 472608
rect 347792 460934 347820 472602
rect 345124 460906 345888 460934
rect 346504 460906 347360 460934
rect 347792 460906 348096 460934
rect 339592 448112 339644 448118
rect 339592 448054 339644 448060
rect 335176 446684 335228 446690
rect 335176 446626 335228 446632
rect 333980 446616 334032 446622
rect 333980 446558 334032 446564
rect 333992 445058 334020 446558
rect 334440 445120 334492 445126
rect 334440 445062 334492 445068
rect 333980 445052 334032 445058
rect 333980 444994 334032 445000
rect 333704 443556 333756 443562
rect 333704 443498 333756 443504
rect 332612 443278 332994 443306
rect 333716 443292 333744 443498
rect 334452 443292 334480 445062
rect 335188 443292 335216 446626
rect 337384 446616 337436 446622
rect 337384 446558 337436 446564
rect 335912 446004 335964 446010
rect 335912 445946 335964 445952
rect 335924 443292 335952 445946
rect 336648 445188 336700 445194
rect 336648 445130 336700 445136
rect 336660 443292 336688 445130
rect 337396 443292 337424 446558
rect 338856 444984 338908 444990
rect 338856 444926 338908 444932
rect 338212 443488 338264 443494
rect 338212 443430 338264 443436
rect 338224 443306 338252 443430
rect 338146 443278 338252 443306
rect 338868 443292 338896 444926
rect 339604 443292 339632 448054
rect 341800 447976 341852 447982
rect 341800 447918 341852 447924
rect 341064 444712 341116 444718
rect 341064 444654 341116 444660
rect 340064 443290 340354 443306
rect 341076 443292 341104 444654
rect 341812 443292 341840 447918
rect 344008 447908 344060 447914
rect 344008 447850 344060 447856
rect 342536 446072 342588 446078
rect 342536 446014 342588 446020
rect 342548 443292 342576 446014
rect 343272 444644 343324 444650
rect 343272 444586 343324 444592
rect 343284 443292 343312 444586
rect 344020 443292 344048 447850
rect 344744 445936 344796 445942
rect 344744 445878 344796 445884
rect 344756 443292 344784 445878
rect 345480 444576 345532 444582
rect 345480 444518 345532 444524
rect 345492 443292 345520 444518
rect 345860 443306 345888 460906
rect 346952 445800 347004 445806
rect 346952 445742 347004 445748
rect 340052 443284 340354 443290
rect 340104 443278 340354 443284
rect 345860 443278 346242 443306
rect 346964 443292 346992 445742
rect 347332 443306 347360 460906
rect 348068 443306 348096 460906
rect 349160 460216 349212 460222
rect 349160 460158 349212 460164
rect 347332 443278 347714 443306
rect 348068 443278 348450 443306
rect 349172 443292 349200 460158
rect 349528 457496 349580 457502
rect 349528 457438 349580 457444
rect 349540 443306 349568 457438
rect 350632 447840 350684 447846
rect 350632 447782 350684 447788
rect 349540 443278 349922 443306
rect 350644 443292 350672 447782
rect 357452 446622 357480 700266
rect 357440 446616 357492 446622
rect 357440 446558 357492 446564
rect 357544 446554 357572 700334
rect 357532 446548 357584 446554
rect 357532 446490 357584 446496
rect 357636 446486 357664 700402
rect 357728 478310 357756 700538
rect 358820 700528 358872 700534
rect 358820 700470 358872 700476
rect 357716 478304 357768 478310
rect 357716 478246 357768 478252
rect 358832 446690 358860 700470
rect 363604 616888 363656 616894
rect 363604 616830 363656 616836
rect 359464 576904 359516 576910
rect 359464 576846 359516 576852
rect 359476 467226 359504 576846
rect 360844 563100 360896 563106
rect 360844 563042 360896 563048
rect 359464 467220 359516 467226
rect 359464 467162 359516 467168
rect 360856 450566 360884 563042
rect 363616 451926 363644 616830
rect 364352 460290 364380 702406
rect 397472 700330 397500 703520
rect 374644 700324 374696 700330
rect 374644 700266 374696 700272
rect 397460 700324 397512 700330
rect 397460 700266 397512 700272
rect 371884 670744 371936 670750
rect 371884 670686 371936 670692
rect 367744 630692 367796 630698
rect 367744 630634 367796 630640
rect 367756 469946 367784 630634
rect 369124 590708 369176 590714
rect 369124 590650 369176 590656
rect 367744 469940 367796 469946
rect 367744 469882 367796 469888
rect 369136 461650 369164 590650
rect 369124 461644 369176 461650
rect 369124 461586 369176 461592
rect 364340 460284 364392 460290
rect 364340 460226 364392 460232
rect 371896 454714 371924 670686
rect 373264 643136 373316 643142
rect 373264 643078 373316 643084
rect 373276 464370 373304 643078
rect 374656 472734 374684 700266
rect 387064 696992 387116 696998
rect 387064 696934 387116 696940
rect 374644 472728 374696 472734
rect 374644 472670 374696 472676
rect 387076 465730 387104 696934
rect 387064 465724 387116 465730
rect 387064 465666 387116 465672
rect 373264 464364 373316 464370
rect 373264 464306 373316 464312
rect 371884 454708 371936 454714
rect 371884 454650 371936 454656
rect 363604 451920 363656 451926
rect 363604 451862 363656 451868
rect 360844 450560 360896 450566
rect 360844 450502 360896 450508
rect 412652 449682 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 429856 699718 429884 703520
rect 462332 700330 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 431224 700324 431276 700330
rect 431224 700266 431276 700272
rect 462320 700324 462372 700330
rect 462320 700266 462372 700272
rect 462964 700324 463016 700330
rect 462964 700266 463016 700272
rect 428464 699712 428516 699718
rect 428464 699654 428516 699660
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 428476 457570 428504 699654
rect 431236 463010 431264 700266
rect 431224 463004 431276 463010
rect 431224 462946 431276 462952
rect 428464 457564 428516 457570
rect 428464 457506 428516 457512
rect 462976 453354 463004 700266
rect 462964 453348 463016 453354
rect 462964 453290 463016 453296
rect 412640 449676 412692 449682
rect 412640 449618 412692 449624
rect 477512 449546 477540 702406
rect 480904 484424 480956 484430
rect 480904 484366 480956 484372
rect 480916 458862 480944 484366
rect 480904 458856 480956 458862
rect 480904 458798 480956 458804
rect 494072 456142 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 496084 536852 496136 536858
rect 496084 536794 496136 536800
rect 496096 468518 496124 536794
rect 496084 468512 496136 468518
rect 496084 468454 496136 468460
rect 494060 456136 494112 456142
rect 494060 456078 494112 456084
rect 477500 449540 477552 449546
rect 477500 449482 477552 449488
rect 527192 448050 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 542372 475386 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 683904 580318 683913
rect 580262 683839 580318 683848
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 580000 630698 580028 630799
rect 579988 630692 580040 630698
rect 579988 630634 580040 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579894 537840 579950 537849
rect 579894 537775 579950 537784
rect 579908 536858 579936 537775
rect 579896 536852 579948 536858
rect 579896 536794 579948 536800
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 542360 475380 542412 475386
rect 542360 475322 542412 475328
rect 580276 471374 580304 683839
rect 580264 471368 580316 471374
rect 580264 471310 580316 471316
rect 527180 448044 527232 448050
rect 527180 447986 527232 447992
rect 358820 446684 358872 446690
rect 358820 446626 358872 446632
rect 357624 446480 357676 446486
rect 357624 446422 357676 446428
rect 362224 446412 362276 446418
rect 362224 446354 362276 446360
rect 360844 446276 360896 446282
rect 360844 446218 360896 446224
rect 359464 446208 359516 446214
rect 359464 446150 359516 446156
rect 356518 445768 356574 445777
rect 356518 445703 356574 445712
rect 351368 444916 351420 444922
rect 351368 444858 351420 444864
rect 351380 443292 351408 444858
rect 352840 444848 352892 444854
rect 352840 444790 352892 444796
rect 351920 443420 351972 443426
rect 351920 443362 351972 443368
rect 351932 443306 351960 443362
rect 351932 443278 352130 443306
rect 352852 443292 352880 444790
rect 355048 444508 355100 444514
rect 355048 444450 355100 444456
rect 355060 443292 355088 444450
rect 356532 443292 356560 445703
rect 340052 443226 340104 443232
rect 353300 443216 353352 443222
rect 353352 443164 353602 443170
rect 353300 443158 353602 443164
rect 353312 443142 353602 443158
rect 355520 443154 355810 443170
rect 355508 443148 355810 443154
rect 355560 443142 355810 443148
rect 355508 443090 355560 443096
rect 354036 443080 354088 443086
rect 354088 443028 354338 443034
rect 354036 443022 354338 443028
rect 354048 443006 354338 443022
rect 356992 443018 357282 443034
rect 356980 443012 357282 443018
rect 357032 443006 357282 443012
rect 356980 442954 357032 442960
rect 359476 442270 359504 446150
rect 359464 442264 359516 442270
rect 359464 442206 359516 442212
rect 230940 440904 230992 440910
rect 230940 440846 230992 440852
rect 230020 398812 230072 398818
rect 230020 398754 230072 398760
rect 229928 372564 229980 372570
rect 229928 372506 229980 372512
rect 229836 346384 229888 346390
rect 229836 346326 229888 346332
rect 238772 310406 240074 310434
rect 238024 309052 238076 309058
rect 238024 308994 238076 309000
rect 229744 244928 229796 244934
rect 229744 244870 229796 244876
rect 237380 174548 237432 174554
rect 237380 174490 237432 174496
rect 158534 159896 158590 159905
rect 158534 159831 158590 159840
rect 165986 159896 166042 159905
rect 165986 159831 166042 159840
rect 173438 159896 173494 159905
rect 173438 159831 173494 159840
rect 156050 159624 156106 159633
rect 156050 159559 156106 159568
rect 156064 159050 156092 159559
rect 156052 159044 156104 159050
rect 156052 158986 156104 158992
rect 158548 158982 158576 159831
rect 166000 159118 166028 159831
rect 173452 159390 173480 159831
rect 206006 159624 206062 159633
rect 206006 159559 206062 159568
rect 173440 159384 173492 159390
rect 173440 159326 173492 159332
rect 206020 159186 206048 159559
rect 231858 159488 231914 159497
rect 231858 159423 231914 159432
rect 213918 159352 213974 159361
rect 213918 159287 213974 159296
rect 206008 159180 206060 159186
rect 206008 159122 206060 159128
rect 165988 159112 166040 159118
rect 165988 159054 166040 159060
rect 158536 158976 158588 158982
rect 158536 158918 158588 158924
rect 168288 158840 168340 158846
rect 168288 158782 168340 158788
rect 160928 158772 160980 158778
rect 160928 158714 160980 158720
rect 120632 158704 120684 158710
rect 116490 158672 116546 158681
rect 116490 158607 116546 158616
rect 117226 158672 117282 158681
rect 119710 158672 119766 158681
rect 117282 158630 117360 158658
rect 117226 158607 117282 158616
rect 116504 157146 116532 158607
rect 117332 157214 117360 158630
rect 119710 158607 119766 158616
rect 120630 158672 120632 158681
rect 160940 158681 160968 158714
rect 168300 158681 168328 158782
rect 120684 158672 120686 158681
rect 120630 158607 120686 158616
rect 121918 158672 121974 158681
rect 121918 158607 121974 158616
rect 123206 158672 123262 158681
rect 123206 158607 123262 158616
rect 126518 158672 126574 158681
rect 126518 158607 126574 158616
rect 128174 158672 128230 158681
rect 128174 158607 128230 158616
rect 128726 158672 128782 158681
rect 128726 158607 128782 158616
rect 130566 158672 130622 158681
rect 130566 158607 130622 158616
rect 131486 158672 131542 158681
rect 131486 158607 131542 158616
rect 132406 158672 132462 158681
rect 132406 158607 132462 158616
rect 133510 158672 133566 158681
rect 133510 158607 133566 158616
rect 134890 158672 134946 158681
rect 134890 158607 134946 158616
rect 158534 158672 158590 158681
rect 158534 158607 158590 158616
rect 159914 158672 159970 158681
rect 159914 158607 159970 158616
rect 160926 158672 160982 158681
rect 160926 158607 160982 158616
rect 168286 158672 168342 158681
rect 168286 158607 168342 158616
rect 119724 158574 119752 158607
rect 119712 158568 119764 158574
rect 119712 158510 119764 158516
rect 118238 158400 118294 158409
rect 118238 158335 118294 158344
rect 117320 157208 117372 157214
rect 117320 157150 117372 157156
rect 116492 157140 116544 157146
rect 116492 157082 116544 157088
rect 118252 156738 118280 158335
rect 121932 157622 121960 158607
rect 121920 157616 121972 157622
rect 121920 157558 121972 157564
rect 123220 157350 123248 158607
rect 126532 158438 126560 158607
rect 126520 158432 126572 158438
rect 126520 158374 126572 158380
rect 128188 158234 128216 158607
rect 128176 158228 128228 158234
rect 128176 158170 128228 158176
rect 128740 158166 128768 158607
rect 130580 158302 130608 158607
rect 130568 158296 130620 158302
rect 130568 158238 130620 158244
rect 128728 158160 128780 158166
rect 128728 158102 128780 158108
rect 131500 158098 131528 158607
rect 131488 158092 131540 158098
rect 131488 158034 131540 158040
rect 132420 158030 132448 158607
rect 133524 158370 133552 158607
rect 133512 158364 133564 158370
rect 133512 158306 133564 158312
rect 133694 158128 133750 158137
rect 133694 158063 133750 158072
rect 132408 158024 132460 158030
rect 132408 157966 132460 157972
rect 124586 157584 124642 157593
rect 124586 157519 124642 157528
rect 123208 157344 123260 157350
rect 123208 157286 123260 157292
rect 118240 156732 118292 156738
rect 118240 156674 118292 156680
rect 124600 154970 124628 157519
rect 125414 157448 125470 157457
rect 125414 157383 125470 157392
rect 124588 154964 124640 154970
rect 124588 154906 124640 154912
rect 125428 154562 125456 157383
rect 133708 155961 133736 158063
rect 134904 157078 134932 158607
rect 135902 158536 135958 158545
rect 135902 158471 135958 158480
rect 137006 158536 137062 158545
rect 137006 158471 137062 158480
rect 138110 158536 138166 158545
rect 138110 158471 138166 158480
rect 148874 158536 148930 158545
rect 148874 158471 148930 158480
rect 134892 157072 134944 157078
rect 134892 157014 134944 157020
rect 135916 157010 135944 158471
rect 136086 157856 136142 157865
rect 136086 157791 136142 157800
rect 135904 157004 135956 157010
rect 135904 156946 135956 156952
rect 133694 155952 133750 155961
rect 133694 155887 133750 155896
rect 136100 155378 136128 157791
rect 137020 156874 137048 158471
rect 138124 156942 138152 158471
rect 141422 158264 141478 158273
rect 141422 158199 141478 158208
rect 141790 158264 141846 158273
rect 141790 158199 141846 158208
rect 144090 158264 144146 158273
rect 144090 158199 144146 158208
rect 146022 158264 146078 158273
rect 146022 158199 146078 158208
rect 146390 158264 146446 158273
rect 146390 158199 146446 158208
rect 140686 157992 140742 158001
rect 140686 157927 140742 157936
rect 140502 157856 140558 157865
rect 140502 157791 140558 157800
rect 138112 156936 138164 156942
rect 138112 156878 138164 156884
rect 137008 156868 137060 156874
rect 137008 156810 137060 156816
rect 140516 155650 140544 157791
rect 140700 155854 140728 157927
rect 140688 155848 140740 155854
rect 140688 155790 140740 155796
rect 140504 155644 140556 155650
rect 140504 155586 140556 155592
rect 136088 155372 136140 155378
rect 136088 155314 136140 155320
rect 125416 154556 125468 154562
rect 125416 154498 125468 154504
rect 141436 153202 141464 158199
rect 141804 155582 141832 158199
rect 143078 157584 143134 157593
rect 143078 157519 143134 157528
rect 141792 155576 141844 155582
rect 141792 155518 141844 155524
rect 143092 154902 143120 157519
rect 144104 156398 144132 158199
rect 145286 157856 145342 157865
rect 145286 157791 145342 157800
rect 144366 157448 144422 157457
rect 144366 157383 144422 157392
rect 144092 156392 144144 156398
rect 144092 156334 144144 156340
rect 143080 154896 143132 154902
rect 143080 154838 143132 154844
rect 141424 153196 141476 153202
rect 141424 153138 141476 153144
rect 144380 153134 144408 157383
rect 144918 156632 144974 156641
rect 144918 156567 144974 156576
rect 144368 153128 144420 153134
rect 144368 153070 144420 153076
rect 135260 152516 135312 152522
rect 135260 152458 135312 152464
rect 121460 149728 121512 149734
rect 121460 149670 121512 149676
rect 115940 141432 115992 141438
rect 115940 141374 115992 141380
rect 107660 140072 107712 140078
rect 107660 140014 107712 140020
rect 103520 137284 103572 137290
rect 103520 137226 103572 137232
rect 102140 93152 102192 93158
rect 102140 93094 102192 93100
rect 99380 89004 99432 89010
rect 99380 88946 99432 88952
rect 99392 16574 99420 88946
rect 93872 16546 94728 16574
rect 95252 16546 95832 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93952 3664 94004 3670
rect 93952 3606 94004 3612
rect 93964 480 93992 3606
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97448 4956 97500 4962
rect 97448 4898 97500 4904
rect 97460 480 97488 4898
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 102152 6914 102180 93094
rect 102232 24132 102284 24138
rect 102232 24074 102284 24080
rect 102244 16574 102272 24074
rect 103532 16574 103560 137226
rect 106280 104168 106332 104174
rect 106280 104110 106332 104116
rect 106292 16574 106320 104110
rect 107672 16574 107700 140014
rect 110420 138712 110472 138718
rect 110420 138654 110472 138660
rect 102244 16546 103376 16574
rect 103532 16546 104112 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 102152 6886 102272 6914
rect 101036 6384 101088 6390
rect 101036 6326 101088 6332
rect 101048 480 101076 6326
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105728 11756 105780 11762
rect 105728 11698 105780 11704
rect 105740 480 105768 11698
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 109040 13116 109092 13122
rect 109040 13058 109092 13064
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 13058
rect 110432 3398 110460 138654
rect 114560 95940 114612 95946
rect 114560 95882 114612 95888
rect 111800 91792 111852 91798
rect 111800 91734 111852 91740
rect 110512 25560 110564 25566
rect 110512 25502 110564 25508
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 25502
rect 111812 16574 111840 91734
rect 113180 26920 113232 26926
rect 113180 26862 113232 26868
rect 113192 16574 113220 26862
rect 114572 16574 114600 95882
rect 115952 16574 115980 141374
rect 120080 130416 120132 130422
rect 120080 130358 120132 130364
rect 118700 127628 118752 127634
rect 118700 127570 118752 127576
rect 117320 86284 117372 86290
rect 117320 86226 117372 86232
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 86226
rect 118712 16574 118740 127570
rect 120092 16574 120120 130358
rect 121472 16574 121500 149670
rect 128360 148368 128412 148374
rect 128360 148310 128412 148316
rect 126980 141500 127032 141506
rect 126980 141442 127032 141448
rect 124220 105596 124272 105602
rect 124220 105538 124272 105544
rect 122840 90364 122892 90370
rect 122840 90306 122892 90312
rect 122852 16574 122880 90306
rect 124232 16574 124260 105538
rect 118712 16546 118832 16574
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 118804 480 118832 16546
rect 119896 14476 119948 14482
rect 119896 14418 119948 14424
rect 119908 480 119936 14418
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 125876 3732 125928 3738
rect 125876 3674 125928 3680
rect 125888 480 125916 3674
rect 126992 480 127020 141442
rect 127072 116612 127124 116618
rect 127072 116554 127124 116560
rect 127084 16574 127112 116554
rect 128372 16574 128400 148310
rect 133880 145580 133932 145586
rect 133880 145522 133932 145528
rect 132500 144220 132552 144226
rect 132500 144162 132552 144168
rect 129740 129056 129792 129062
rect 129740 128998 129792 129004
rect 129752 16574 129780 128998
rect 131120 108316 131172 108322
rect 131120 108258 131172 108264
rect 131132 16574 131160 108258
rect 132512 16574 132540 144162
rect 127084 16546 128216 16574
rect 128372 16546 128952 16574
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 132512 16546 133000 16574
rect 128188 480 128216 16546
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 130580 480 130608 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 132972 480 133000 16546
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 133892 354 133920 145522
rect 135272 3806 135300 152458
rect 139400 146940 139452 146946
rect 139400 146882 139452 146888
rect 136640 123480 136692 123486
rect 136640 123422 136692 123428
rect 135352 102808 135404 102814
rect 135352 102750 135404 102756
rect 135260 3800 135312 3806
rect 135260 3742 135312 3748
rect 135364 3482 135392 102750
rect 136652 16574 136680 123422
rect 138020 101448 138072 101454
rect 138020 101390 138072 101396
rect 138032 16574 138060 101390
rect 139412 16574 139440 146882
rect 143540 142860 143592 142866
rect 143540 142802 143592 142808
rect 140780 122120 140832 122126
rect 140780 122062 140832 122068
rect 140792 16574 140820 122062
rect 142160 19984 142212 19990
rect 142160 19926 142212 19932
rect 136652 16546 137232 16574
rect 138032 16546 138888 16574
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 136456 3800 136508 3806
rect 136456 3742 136508 3748
rect 135272 3454 135392 3482
rect 135272 480 135300 3454
rect 136468 480 136496 3742
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 138860 480 138888 16546
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142172 354 142200 19926
rect 143552 480 143580 142802
rect 143632 134564 143684 134570
rect 143632 134506 143684 134512
rect 143644 16574 143672 134506
rect 144932 16574 144960 156567
rect 145300 155514 145328 157791
rect 145288 155508 145340 155514
rect 145288 155450 145340 155456
rect 146036 153066 146064 158199
rect 146404 155446 146432 158199
rect 147678 157856 147734 157865
rect 147678 157791 147734 157800
rect 146392 155440 146444 155446
rect 146392 155382 146444 155388
rect 147692 155310 147720 157791
rect 148506 157448 148562 157457
rect 148506 157383 148562 157392
rect 147680 155304 147732 155310
rect 147680 155246 147732 155252
rect 146024 153060 146076 153066
rect 146024 153002 146076 153008
rect 148520 152998 148548 157383
rect 148888 156806 148916 158471
rect 150990 158264 151046 158273
rect 150990 158199 151046 158208
rect 149886 157448 149942 157457
rect 149886 157383 149942 157392
rect 148876 156800 148928 156806
rect 148876 156742 148928 156748
rect 149900 154290 149928 157383
rect 149888 154284 149940 154290
rect 149888 154226 149940 154232
rect 148508 152992 148560 152998
rect 148508 152934 148560 152940
rect 151004 152930 151032 158199
rect 158548 157962 158576 158607
rect 158536 157956 158588 157962
rect 158536 157898 158588 157904
rect 159928 157894 159956 158607
rect 195886 158536 195942 158545
rect 195886 158471 195942 158480
rect 178866 158400 178922 158409
rect 178866 158335 178922 158344
rect 181810 158400 181866 158409
rect 181810 158335 181866 158344
rect 184018 158400 184074 158409
rect 184018 158335 184074 158344
rect 159916 157888 159968 157894
rect 159916 157830 159968 157836
rect 151358 157448 151414 157457
rect 151358 157383 151414 157392
rect 152646 157448 152702 157457
rect 152646 157383 152702 157392
rect 154118 157448 154174 157457
rect 154118 157383 154174 157392
rect 154486 157448 154542 157457
rect 154486 157383 154542 157392
rect 155774 157448 155830 157457
rect 155774 157383 155830 157392
rect 157062 157448 157118 157457
rect 157062 157383 157118 157392
rect 151372 154222 151400 157383
rect 152660 154358 152688 157383
rect 153198 155272 153254 155281
rect 153198 155207 153254 155216
rect 152648 154352 152700 154358
rect 152648 154294 152700 154300
rect 151360 154216 151412 154222
rect 151360 154158 151412 154164
rect 150992 152924 151044 152930
rect 150992 152866 151044 152872
rect 146300 151088 146352 151094
rect 146300 151030 146352 151036
rect 146312 16574 146340 151030
rect 150440 145648 150492 145654
rect 150440 145590 150492 145596
rect 147680 120760 147732 120766
rect 147680 120702 147732 120708
rect 147692 16574 147720 120702
rect 149060 100020 149112 100026
rect 149060 99962 149112 99968
rect 149072 16574 149100 99962
rect 150452 16574 150480 145590
rect 151820 133204 151872 133210
rect 151820 133146 151872 133152
rect 143644 16546 144776 16574
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 150452 16546 150664 16574
rect 144748 480 144776 16546
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150636 480 150664 16546
rect 151832 480 151860 133146
rect 151912 98660 151964 98666
rect 151912 98602 151964 98608
rect 151924 16574 151952 98602
rect 153212 16574 153240 155207
rect 154132 154494 154160 157383
rect 154120 154488 154172 154494
rect 154120 154430 154172 154436
rect 154500 153814 154528 157383
rect 155788 154426 155816 157383
rect 157076 154834 157104 157383
rect 175278 156768 175334 156777
rect 175278 156703 175334 156712
rect 157064 154828 157116 154834
rect 157064 154770 157116 154776
rect 155776 154420 155828 154426
rect 155776 154362 155828 154368
rect 168380 153876 168432 153882
rect 168380 153818 168432 153824
rect 154488 153808 154540 153814
rect 154488 153750 154540 153756
rect 157340 149796 157392 149802
rect 157340 149738 157392 149744
rect 155960 135924 156012 135930
rect 155960 135866 156012 135872
rect 154580 119400 154632 119406
rect 154580 119342 154632 119348
rect 154592 16574 154620 119342
rect 155972 16574 156000 135866
rect 157352 16574 157380 149738
rect 161480 140140 161532 140146
rect 161480 140082 161532 140088
rect 158720 117972 158772 117978
rect 158720 117914 158772 117920
rect 158732 16574 158760 117914
rect 160100 21412 160152 21418
rect 160100 21354 160152 21360
rect 151924 16546 153056 16574
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 153028 480 153056 16546
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 480 160140 21354
rect 161492 16574 161520 140082
rect 165620 138780 165672 138786
rect 165620 138722 165672 138728
rect 162860 115252 162912 115258
rect 162860 115194 162912 115200
rect 162872 16574 162900 115194
rect 165632 16574 165660 138722
rect 167000 113824 167052 113830
rect 167000 113766 167052 113772
rect 167012 16574 167040 113766
rect 161492 16546 162072 16574
rect 162872 16546 163728 16574
rect 165632 16546 166120 16574
rect 167012 16546 167224 16574
rect 161296 3800 161348 3806
rect 161296 3742 161348 3748
rect 161308 480 161336 3742
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163700 480 163728 16546
rect 164884 5024 164936 5030
rect 164884 4966 164936 4972
rect 164896 480 164924 4966
rect 166092 480 166120 16546
rect 167196 480 167224 16546
rect 168392 480 168420 153818
rect 169760 124908 169812 124914
rect 169760 124850 169812 124856
rect 169772 16574 169800 124850
rect 173900 112464 173952 112470
rect 173900 112406 173952 112412
rect 169772 16546 170352 16574
rect 169576 5092 169628 5098
rect 169576 5034 169628 5040
rect 169588 480 169616 5034
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 173164 6452 173216 6458
rect 173164 6394 173216 6400
rect 171968 3868 172020 3874
rect 171968 3810 172020 3816
rect 171980 480 172008 3810
rect 173176 480 173204 6394
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 173912 354 173940 112406
rect 175292 16574 175320 156703
rect 178880 156670 178908 158335
rect 178868 156664 178920 156670
rect 178868 156606 178920 156612
rect 181824 156602 181852 158335
rect 181812 156596 181864 156602
rect 181812 156538 181864 156544
rect 184032 156534 184060 158335
rect 185950 158264 186006 158273
rect 185950 158199 186006 158208
rect 184020 156528 184072 156534
rect 184020 156470 184072 156476
rect 185964 156466 185992 158199
rect 185952 156460 186004 156466
rect 185952 156402 186004 156408
rect 178038 155408 178094 155417
rect 178038 155343 178094 155352
rect 178052 16574 178080 155343
rect 195900 155242 195928 158471
rect 198462 157584 198518 157593
rect 198462 157519 198518 157528
rect 201038 157584 201094 157593
rect 201038 157519 201094 157528
rect 203430 157584 203486 157593
rect 203430 157519 203486 157528
rect 195888 155236 195940 155242
rect 195888 155178 195940 155184
rect 198476 155174 198504 157519
rect 198464 155168 198516 155174
rect 198464 155110 198516 155116
rect 201052 155106 201080 157519
rect 202878 156904 202934 156913
rect 202878 156839 202934 156848
rect 201040 155100 201092 155106
rect 201040 155042 201092 155048
rect 193220 153944 193272 153950
rect 193220 153886 193272 153892
rect 182180 151156 182232 151162
rect 182180 151098 182232 151104
rect 179420 134632 179472 134638
rect 179420 134574 179472 134580
rect 179432 16574 179460 134574
rect 180800 126268 180852 126274
rect 180800 126210 180852 126216
rect 180812 16574 180840 126210
rect 175292 16546 175504 16574
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 175476 480 175504 16546
rect 177856 7676 177908 7682
rect 177856 7618 177908 7624
rect 176660 6520 176712 6526
rect 176660 6462 176712 6468
rect 176672 480 176700 6462
rect 177868 480 177896 7618
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182192 354 182220 151098
rect 184940 149864 184992 149870
rect 184940 149806 184992 149812
rect 183560 133272 183612 133278
rect 183560 133214 183612 133220
rect 183572 16574 183600 133214
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 184952 11830 184980 149806
rect 186320 144288 186372 144294
rect 186320 144230 186372 144236
rect 185032 111104 185084 111110
rect 185032 111046 185084 111052
rect 184940 11824 184992 11830
rect 184940 11766 184992 11772
rect 185044 6914 185072 111046
rect 186332 16574 186360 144230
rect 187700 131844 187752 131850
rect 187700 131786 187752 131792
rect 187712 16574 187740 131786
rect 190460 131776 190512 131782
rect 190460 131718 190512 131724
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 186136 11824 186188 11830
rect 186136 11766 186188 11772
rect 184952 6886 185072 6914
rect 184952 480 184980 6886
rect 186148 480 186176 11766
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 189724 5160 189776 5166
rect 189724 5102 189776 5108
rect 189736 480 189764 5102
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 354 190500 131718
rect 191840 109744 191892 109750
rect 191840 109686 191892 109692
rect 191852 16574 191880 109686
rect 191852 16546 192064 16574
rect 192036 480 192064 16546
rect 193232 480 193260 153886
rect 195978 152416 196034 152425
rect 195978 152351 196034 152360
rect 193312 130484 193364 130490
rect 193312 130426 193364 130432
rect 193324 16574 193352 130426
rect 194600 17264 194652 17270
rect 194600 17206 194652 17212
rect 194612 16574 194640 17206
rect 195992 16574 196020 152351
rect 200120 147008 200172 147014
rect 200120 146950 200172 146956
rect 197360 142928 197412 142934
rect 197360 142870 197412 142876
rect 197372 16574 197400 142870
rect 198740 129124 198792 129130
rect 198740 129066 198792 129072
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 195992 16546 196848 16574
rect 197372 16546 197952 16574
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196820 480 196848 16546
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 129066
rect 200132 16574 200160 146950
rect 201500 141568 201552 141574
rect 201500 141510 201552 141516
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 480 201540 141510
rect 201592 106956 201644 106962
rect 201592 106898 201644 106904
rect 201604 16574 201632 106898
rect 202892 16574 202920 156839
rect 203444 155038 203472 157519
rect 203432 155032 203484 155038
rect 203432 154974 203484 154980
rect 208400 154012 208452 154018
rect 208400 153954 208452 153960
rect 205640 130552 205692 130558
rect 205640 130494 205692 130500
rect 204260 127696 204312 127702
rect 204260 127638 204312 127644
rect 204272 16574 204300 127638
rect 205652 16574 205680 130494
rect 208412 16574 208440 153954
rect 209780 142996 209832 143002
rect 209780 142938 209832 142944
rect 201604 16546 202736 16574
rect 202892 16546 203472 16574
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 208412 16546 208624 16574
rect 202708 480 202736 16546
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203444 354 203472 16546
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 207388 5228 207440 5234
rect 207388 5170 207440 5176
rect 207400 480 207428 5170
rect 208596 480 208624 16546
rect 209792 480 209820 142938
rect 211160 140208 211212 140214
rect 211160 140150 211212 140156
rect 211172 16574 211200 140150
rect 212540 18624 212592 18630
rect 212540 18566 212592 18572
rect 212552 16574 212580 18566
rect 213932 16574 213960 159287
rect 220818 155544 220874 155553
rect 220818 155479 220874 155488
rect 218060 145716 218112 145722
rect 218060 145658 218112 145664
rect 216680 144356 216732 144362
rect 216680 144298 216732 144304
rect 215298 138680 215354 138689
rect 215298 138615 215354 138624
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 213932 16546 214512 16574
rect 210976 5296 211028 5302
rect 210976 5238 211028 5244
rect 210988 480 211016 5238
rect 203862 354 203974 480
rect 203444 326 203974 354
rect 203862 -960 203974 326
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 138615
rect 216692 16574 216720 144298
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 480 218100 145658
rect 218152 126336 218204 126342
rect 218152 126278 218204 126284
rect 218164 16574 218192 126278
rect 219440 105664 219492 105670
rect 219440 105606 219492 105612
rect 219452 16574 219480 105606
rect 220832 16574 220860 155479
rect 227720 154080 227772 154086
rect 227720 154022 227772 154028
rect 224960 148436 225012 148442
rect 224960 148378 225012 148384
rect 222198 146976 222254 146985
rect 222198 146911 222254 146920
rect 222212 16574 222240 146911
rect 223578 127664 223634 127673
rect 223578 127599 223634 127608
rect 218164 16546 219296 16574
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 127599
rect 224972 16574 225000 148378
rect 226340 137352 226392 137358
rect 226340 137294 226392 137300
rect 224972 16546 225184 16574
rect 225156 480 225184 16546
rect 226352 480 226380 137294
rect 227732 16574 227760 154022
rect 229100 124976 229152 124982
rect 229100 124918 229152 124924
rect 229112 16574 229140 124918
rect 230480 104236 230532 104242
rect 230480 104178 230532 104184
rect 230492 16574 230520 104178
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 227536 10396 227588 10402
rect 227536 10338 227588 10344
rect 227548 480 227576 10338
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 159423
rect 234620 157820 234672 157826
rect 234620 157762 234672 157768
rect 234632 156738 234660 157762
rect 234620 156732 234672 156738
rect 234620 156674 234672 156680
rect 236000 89140 236052 89146
rect 236000 89082 236052 89088
rect 233240 89072 233292 89078
rect 233240 89014 233292 89020
rect 233252 16574 233280 89014
rect 236012 16574 236040 89082
rect 237392 16574 237420 174490
rect 238036 86290 238064 308994
rect 238208 308984 238260 308990
rect 238208 308926 238260 308932
rect 238116 174684 238168 174690
rect 238116 174626 238168 174632
rect 238024 86284 238076 86290
rect 238024 86226 238076 86232
rect 233252 16546 233464 16574
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 233436 480 233464 16546
rect 234620 6656 234672 6662
rect 234620 6598 234672 6604
rect 234632 480 234660 6598
rect 235816 6588 235868 6594
rect 235816 6530 235868 6536
rect 235828 480 235856 6530
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 238128 3738 238156 174626
rect 238220 159118 238248 308926
rect 238300 297628 238352 297634
rect 238300 297570 238352 297576
rect 238208 159112 238260 159118
rect 238208 159054 238260 159060
rect 238312 158137 238340 297570
rect 238484 254584 238536 254590
rect 238484 254526 238536 254532
rect 238392 170400 238444 170406
rect 238392 170342 238444 170348
rect 238404 159594 238432 170342
rect 238392 159588 238444 159594
rect 238392 159530 238444 159536
rect 238298 158128 238354 158137
rect 238298 158063 238354 158072
rect 238496 158001 238524 254526
rect 238576 167680 238628 167686
rect 238576 167622 238628 167628
rect 238588 159662 238616 167622
rect 238576 159656 238628 159662
rect 238576 159598 238628 159604
rect 238482 157992 238538 158001
rect 238482 157927 238538 157936
rect 238772 94518 238800 310406
rect 240244 308496 240272 310420
rect 240152 308468 240272 308496
rect 240152 307086 240180 308468
rect 240428 308394 240456 310420
rect 240244 308366 240456 308394
rect 240140 307080 240192 307086
rect 240140 307022 240192 307028
rect 240244 304298 240272 308366
rect 240612 308292 240640 310420
rect 240796 308446 240824 310420
rect 240784 308440 240836 308446
rect 240784 308382 240836 308388
rect 240336 308264 240640 308292
rect 240232 304292 240284 304298
rect 240232 304234 240284 304240
rect 240336 280838 240364 308264
rect 240980 308122 241008 310420
rect 240428 308094 241008 308122
rect 240324 280832 240376 280838
rect 240324 280774 240376 280780
rect 240428 265674 240456 308094
rect 240508 308032 240560 308038
rect 240508 307974 240560 307980
rect 240520 279478 240548 307974
rect 241164 302938 241192 310420
rect 241348 308038 241376 310420
rect 241532 308394 241560 310420
rect 241716 308718 241744 310420
rect 241704 308712 241756 308718
rect 241704 308654 241756 308660
rect 241900 308496 241928 310420
rect 241808 308468 241928 308496
rect 241532 308366 241744 308394
rect 241612 308304 241664 308310
rect 241612 308246 241664 308252
rect 241336 308032 241388 308038
rect 241336 307974 241388 307980
rect 241624 304366 241652 308246
rect 241612 304360 241664 304366
rect 241612 304302 241664 304308
rect 241152 302932 241204 302938
rect 241152 302874 241204 302880
rect 240508 279472 240560 279478
rect 240508 279414 240560 279420
rect 240416 265668 240468 265674
rect 240416 265610 240468 265616
rect 241716 260166 241744 308366
rect 241808 308310 241836 308468
rect 242084 308394 242112 310420
rect 241900 308366 242112 308394
rect 241796 308304 241848 308310
rect 241796 308246 241848 308252
rect 241796 308168 241848 308174
rect 241796 308110 241848 308116
rect 241808 264246 241836 308110
rect 241900 294642 241928 308366
rect 241980 308304 242032 308310
rect 242268 308292 242296 310420
rect 242452 308310 242480 310420
rect 241980 308246 242032 308252
rect 242084 308264 242296 308292
rect 242440 308304 242492 308310
rect 241888 294636 241940 294642
rect 241888 294578 241940 294584
rect 241796 264240 241848 264246
rect 241796 264182 241848 264188
rect 241704 260160 241756 260166
rect 241704 260102 241756 260108
rect 240138 175944 240194 175953
rect 240138 175879 240194 175888
rect 239404 173188 239456 173194
rect 239404 173130 239456 173136
rect 238760 94512 238812 94518
rect 238760 94454 238812 94460
rect 238760 89208 238812 89214
rect 238760 89150 238812 89156
rect 238772 16574 238800 89150
rect 238772 16546 239352 16574
rect 238116 3732 238168 3738
rect 238116 3674 238168 3680
rect 239324 480 239352 16546
rect 239416 3874 239444 173130
rect 239404 3868 239456 3874
rect 239404 3810 239456 3816
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 175879
rect 241612 89276 241664 89282
rect 241612 89218 241664 89224
rect 241624 16574 241652 89218
rect 241624 16546 241744 16574
rect 241716 480 241744 16546
rect 241992 4826 242020 308246
rect 242084 250510 242112 308264
rect 242440 308246 242492 308252
rect 242164 307964 242216 307970
rect 242164 307906 242216 307912
rect 242072 250504 242124 250510
rect 242072 250446 242124 250452
rect 242176 25566 242204 307906
rect 242636 300150 242664 310420
rect 242820 308174 242848 310420
rect 243004 308514 243032 310420
rect 243188 308922 243216 310420
rect 243176 308916 243228 308922
rect 243176 308858 243228 308864
rect 242992 308508 243044 308514
rect 242992 308450 243044 308456
rect 243084 308440 243136 308446
rect 243372 308394 243400 310420
rect 243556 308446 243584 310420
rect 243740 308650 243768 310420
rect 243728 308644 243780 308650
rect 243728 308586 243780 308592
rect 243084 308382 243136 308388
rect 242992 308372 243044 308378
rect 242992 308314 243044 308320
rect 242808 308168 242860 308174
rect 242808 308110 242860 308116
rect 242624 300144 242676 300150
rect 242624 300086 242676 300092
rect 243004 284986 243032 308314
rect 243096 290494 243124 308382
rect 243188 308366 243400 308394
rect 243544 308440 243596 308446
rect 243544 308382 243596 308388
rect 243188 298790 243216 308366
rect 243924 308292 243952 310420
rect 244108 308378 244136 310420
rect 244292 308394 244320 310420
rect 244476 309126 244504 310420
rect 244464 309120 244516 309126
rect 244464 309062 244516 309068
rect 244660 308496 244688 310420
rect 244660 308468 244780 308496
rect 244096 308372 244148 308378
rect 244292 308366 244688 308394
rect 244096 308314 244148 308320
rect 243280 308264 243952 308292
rect 244556 308304 244608 308310
rect 243176 298784 243228 298790
rect 243176 298726 243228 298732
rect 243084 290488 243136 290494
rect 243084 290430 243136 290436
rect 242992 284980 243044 284986
rect 242992 284922 243044 284928
rect 243280 28286 243308 308264
rect 244556 308246 244608 308252
rect 244464 308236 244516 308242
rect 244464 308178 244516 308184
rect 243542 308136 243598 308145
rect 243542 308071 243598 308080
rect 243636 308100 243688 308106
rect 243556 159050 243584 308071
rect 243636 308042 243688 308048
rect 243648 246362 243676 308042
rect 243728 308032 243780 308038
rect 243728 307974 243780 307980
rect 243740 247722 243768 307974
rect 244476 305658 244504 308178
rect 244464 305652 244516 305658
rect 244464 305594 244516 305600
rect 244568 287706 244596 308246
rect 244660 303006 244688 308366
rect 244752 307154 244780 308468
rect 244740 307148 244792 307154
rect 244740 307090 244792 307096
rect 244648 303000 244700 303006
rect 244648 302942 244700 302948
rect 244844 289134 244872 310420
rect 244924 308576 244976 308582
rect 244924 308518 244976 308524
rect 244832 289128 244884 289134
rect 244832 289070 244884 289076
rect 244556 287700 244608 287706
rect 244556 287642 244608 287648
rect 243728 247716 243780 247722
rect 243728 247658 243780 247664
rect 243636 246356 243688 246362
rect 243636 246298 243688 246304
rect 243544 159044 243596 159050
rect 243544 158986 243596 158992
rect 243268 28280 243320 28286
rect 243268 28222 243320 28228
rect 242164 25560 242216 25566
rect 242164 25502 242216 25508
rect 242900 6724 242952 6730
rect 242900 6666 242952 6672
rect 241980 4820 242032 4826
rect 241980 4762 242032 4768
rect 242912 480 242940 6666
rect 244936 6186 244964 308518
rect 245028 308038 245056 310420
rect 245212 308242 245240 310420
rect 245396 308310 245424 310420
rect 245580 308786 245608 310420
rect 245568 308780 245620 308786
rect 245568 308722 245620 308728
rect 245764 308496 245792 310420
rect 245672 308468 245792 308496
rect 245384 308304 245436 308310
rect 245384 308246 245436 308252
rect 245200 308236 245252 308242
rect 245200 308178 245252 308184
rect 245672 308174 245700 308468
rect 245948 308394 245976 310420
rect 246132 308394 246160 310420
rect 246316 308446 246344 310420
rect 245764 308366 245976 308394
rect 246040 308366 246160 308394
rect 246304 308440 246356 308446
rect 246304 308382 246356 308388
rect 245660 308168 245712 308174
rect 245660 308110 245712 308116
rect 245016 308032 245068 308038
rect 245016 307974 245068 307980
rect 245764 301510 245792 308366
rect 245936 308304 245988 308310
rect 245936 308246 245988 308252
rect 245844 308236 245896 308242
rect 245844 308178 245896 308184
rect 245752 301504 245804 301510
rect 245752 301446 245804 301452
rect 245856 282198 245884 308178
rect 245948 283626 245976 308246
rect 245936 283620 245988 283626
rect 245936 283562 245988 283568
rect 245844 282192 245896 282198
rect 245844 282134 245896 282140
rect 245752 174616 245804 174622
rect 245752 174558 245804 174564
rect 245764 16574 245792 174558
rect 245764 16546 245976 16574
rect 244924 6180 244976 6186
rect 244924 6122 244976 6128
rect 245200 4820 245252 4826
rect 245200 4762 245252 4768
rect 244096 3732 244148 3738
rect 244096 3674 244148 3680
rect 244108 480 244136 3674
rect 245212 480 245240 4762
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 246040 7614 246068 308366
rect 246500 308292 246528 310420
rect 246684 308854 246712 310420
rect 246672 308848 246724 308854
rect 246672 308790 246724 308796
rect 246672 308644 246724 308650
rect 246672 308586 246724 308592
rect 246580 308508 246632 308514
rect 246580 308450 246632 308456
rect 246132 308264 246528 308292
rect 246132 262886 246160 308264
rect 246212 308168 246264 308174
rect 246212 308110 246264 308116
rect 246224 297430 246252 308110
rect 246304 307828 246356 307834
rect 246304 307770 246356 307776
rect 246212 297424 246264 297430
rect 246212 297366 246264 297372
rect 246120 262880 246172 262886
rect 246120 262822 246172 262828
rect 246316 22778 246344 307770
rect 246592 296714 246620 308450
rect 246684 307834 246712 308586
rect 246868 308242 246896 310420
rect 247052 308582 247080 310420
rect 247040 308576 247092 308582
rect 247040 308518 247092 308524
rect 247236 308514 247264 310420
rect 247224 308508 247276 308514
rect 247224 308450 247276 308456
rect 247420 308394 247448 310420
rect 247604 308514 247632 310420
rect 247788 308514 247816 310420
rect 247592 308508 247644 308514
rect 247592 308450 247644 308456
rect 247776 308508 247828 308514
rect 247776 308450 247828 308456
rect 247972 308394 248000 310420
rect 248156 308938 248184 310420
rect 248156 308910 248276 308938
rect 248144 308848 248196 308854
rect 248144 308790 248196 308796
rect 248052 308712 248104 308718
rect 248052 308654 248104 308660
rect 247144 308366 247448 308394
rect 247512 308366 248000 308394
rect 246856 308236 246908 308242
rect 246856 308178 246908 308184
rect 246672 307828 246724 307834
rect 246672 307770 246724 307776
rect 246408 296686 246620 296714
rect 246408 87650 246436 296686
rect 246396 87644 246448 87650
rect 246396 87586 246448 87592
rect 246304 22772 246356 22778
rect 246304 22714 246356 22720
rect 246028 7608 246080 7614
rect 246028 7550 246080 7556
rect 247144 3466 247172 308366
rect 247224 308304 247276 308310
rect 247224 308246 247276 308252
rect 247236 4894 247264 308246
rect 247408 308236 247460 308242
rect 247408 308178 247460 308184
rect 247316 308168 247368 308174
rect 247316 308110 247368 308116
rect 247328 6254 247356 308110
rect 247420 286346 247448 308178
rect 247408 286340 247460 286346
rect 247408 286282 247460 286288
rect 247408 22772 247460 22778
rect 247408 22714 247460 22720
rect 247316 6248 247368 6254
rect 247316 6190 247368 6196
rect 247224 4888 247276 4894
rect 247224 4830 247276 4836
rect 247420 3482 247448 22714
rect 247512 16574 247540 308366
rect 247960 308304 248012 308310
rect 247960 308246 248012 308252
rect 247684 307828 247736 307834
rect 247684 307770 247736 307776
rect 247696 24138 247724 307770
rect 247972 307222 248000 308246
rect 247960 307216 248012 307222
rect 247960 307158 248012 307164
rect 248064 296714 248092 308654
rect 248156 307834 248184 308790
rect 248248 308174 248276 308910
rect 248340 308582 248368 310420
rect 248420 308780 248472 308786
rect 248420 308722 248472 308728
rect 248328 308576 248380 308582
rect 248328 308518 248380 308524
rect 248432 308514 248460 308722
rect 248420 308508 248472 308514
rect 248420 308450 248472 308456
rect 248328 308440 248380 308446
rect 248328 308382 248380 308388
rect 248236 308168 248288 308174
rect 248236 308110 248288 308116
rect 248340 307970 248368 308382
rect 248420 308372 248472 308378
rect 248420 308314 248472 308320
rect 248328 307964 248380 307970
rect 248328 307906 248380 307912
rect 248144 307828 248196 307834
rect 248144 307770 248196 307776
rect 247788 296686 248092 296714
rect 247788 89010 247816 296686
rect 248432 296002 248460 308314
rect 248524 298858 248552 310420
rect 248604 308304 248656 308310
rect 248604 308246 248656 308252
rect 248512 298852 248564 298858
rect 248512 298794 248564 298800
rect 248420 295996 248472 296002
rect 248420 295938 248472 295944
rect 248616 273970 248644 308246
rect 248708 275330 248736 310420
rect 248788 308508 248840 308514
rect 248788 308450 248840 308456
rect 248800 297498 248828 308450
rect 248892 308394 248920 310420
rect 249076 308514 249104 310420
rect 249064 308508 249116 308514
rect 249064 308450 249116 308456
rect 248892 308366 249196 308394
rect 248880 308032 248932 308038
rect 248880 307974 248932 307980
rect 248788 297492 248840 297498
rect 248788 297434 248840 297440
rect 248696 275324 248748 275330
rect 248696 275266 248748 275272
rect 248604 273964 248656 273970
rect 248604 273906 248656 273912
rect 248892 253230 248920 307974
rect 249168 296714 249196 308366
rect 249260 308310 249288 310420
rect 249248 308304 249300 308310
rect 249248 308246 249300 308252
rect 249444 308038 249472 310420
rect 249628 308378 249656 310420
rect 249616 308372 249668 308378
rect 249616 308314 249668 308320
rect 249812 308122 249840 310420
rect 249996 308258 250024 310420
rect 249996 308230 250116 308258
rect 249812 308094 250024 308122
rect 249432 308032 249484 308038
rect 249432 307974 249484 307980
rect 249800 308032 249852 308038
rect 249800 307974 249852 307980
rect 249892 308032 249944 308038
rect 249892 307974 249944 307980
rect 249812 307290 249840 307974
rect 249800 307284 249852 307290
rect 249800 307226 249852 307232
rect 249904 300218 249932 307974
rect 249892 300212 249944 300218
rect 249892 300154 249944 300160
rect 248984 296686 249196 296714
rect 248984 258738 249012 296686
rect 249996 272542 250024 308094
rect 250088 285054 250116 308230
rect 250180 308106 250208 310420
rect 250260 308440 250312 308446
rect 250260 308382 250312 308388
rect 250168 308100 250220 308106
rect 250168 308042 250220 308048
rect 250168 307964 250220 307970
rect 250168 307906 250220 307912
rect 250180 294710 250208 307906
rect 250168 294704 250220 294710
rect 250168 294646 250220 294652
rect 250076 285048 250128 285054
rect 250076 284990 250128 284996
rect 249984 272536 250036 272542
rect 249984 272478 250036 272484
rect 248972 258732 249024 258738
rect 248972 258674 249024 258680
rect 248880 253224 248932 253230
rect 248880 253166 248932 253172
rect 247776 89004 247828 89010
rect 247776 88946 247828 88952
rect 247684 24132 247736 24138
rect 247684 24074 247736 24080
rect 247512 16546 247724 16574
rect 247696 3534 247724 16546
rect 250272 6322 250300 308382
rect 250364 271182 250392 310420
rect 250548 308038 250576 310420
rect 250536 308032 250588 308038
rect 250536 307974 250588 307980
rect 250732 307970 250760 310420
rect 250916 308446 250944 310420
rect 250904 308440 250956 308446
rect 250904 308382 250956 308388
rect 250720 307964 250772 307970
rect 250720 307906 250772 307912
rect 251100 298926 251128 310420
rect 251180 308440 251232 308446
rect 251180 308382 251232 308388
rect 251088 298920 251140 298926
rect 251088 298862 251140 298868
rect 251192 291854 251220 308382
rect 251284 305726 251312 310420
rect 251468 308394 251496 310420
rect 251376 308366 251496 308394
rect 251272 305720 251324 305726
rect 251272 305662 251324 305668
rect 251180 291848 251232 291854
rect 251180 291790 251232 291796
rect 250352 271176 250404 271182
rect 250352 271118 250404 271124
rect 251376 269822 251404 308366
rect 251456 308304 251508 308310
rect 251456 308246 251508 308252
rect 251468 283694 251496 308246
rect 251548 306876 251600 306882
rect 251548 306818 251600 306824
rect 251560 290562 251588 306818
rect 251548 290556 251600 290562
rect 251548 290498 251600 290504
rect 251456 283688 251508 283694
rect 251456 283630 251508 283636
rect 251364 269816 251416 269822
rect 251364 269758 251416 269764
rect 251652 251870 251680 310420
rect 251836 308446 251864 310420
rect 251824 308440 251876 308446
rect 251824 308382 251876 308388
rect 252020 296714 252048 310420
rect 252204 308310 252232 310420
rect 252192 308304 252244 308310
rect 252192 308246 252244 308252
rect 252388 306882 252416 310420
rect 252572 308310 252600 310420
rect 252652 308440 252704 308446
rect 252652 308382 252704 308388
rect 252560 308304 252612 308310
rect 252560 308246 252612 308252
rect 252376 306876 252428 306882
rect 252376 306818 252428 306824
rect 252664 303074 252692 308382
rect 252652 303068 252704 303074
rect 252652 303010 252704 303016
rect 251744 296686 252048 296714
rect 251744 268394 251772 296686
rect 252756 282266 252784 310420
rect 252940 308446 252968 310420
rect 252928 308440 252980 308446
rect 253124 308394 253152 310420
rect 252928 308382 252980 308388
rect 252836 308372 252888 308378
rect 252836 308314 252888 308320
rect 253032 308366 253152 308394
rect 252848 289202 252876 308314
rect 252928 308236 252980 308242
rect 252928 308178 252980 308184
rect 252836 289196 252888 289202
rect 252836 289138 252888 289144
rect 252744 282260 252796 282266
rect 252744 282202 252796 282208
rect 251732 268388 251784 268394
rect 251732 268330 251784 268336
rect 251640 251864 251692 251870
rect 251640 251806 251692 251812
rect 252940 8974 252968 308178
rect 253032 265742 253060 308366
rect 253112 308304 253164 308310
rect 253112 308246 253164 308252
rect 253124 296070 253152 308246
rect 253204 308100 253256 308106
rect 253204 308042 253256 308048
rect 253112 296064 253164 296070
rect 253112 296006 253164 296012
rect 253020 265736 253072 265742
rect 253020 265678 253072 265684
rect 253216 14482 253244 308042
rect 253308 305794 253336 310420
rect 253492 308378 253520 310420
rect 253480 308372 253532 308378
rect 253480 308314 253532 308320
rect 253676 308242 253704 310420
rect 253860 308650 253888 310420
rect 253848 308644 253900 308650
rect 253848 308586 253900 308592
rect 253664 308236 253716 308242
rect 253664 308178 253716 308184
rect 253940 307012 253992 307018
rect 253940 306954 253992 306960
rect 253296 305788 253348 305794
rect 253296 305730 253348 305736
rect 253952 304434 253980 306954
rect 254044 306898 254072 310420
rect 254228 307018 254256 310420
rect 254216 307012 254268 307018
rect 254216 306954 254268 306960
rect 254044 306870 254348 306898
rect 254216 306264 254268 306270
rect 254216 306206 254268 306212
rect 253940 304428 253992 304434
rect 253940 304370 253992 304376
rect 254124 304292 254176 304298
rect 254124 304234 254176 304240
rect 253204 14476 253256 14482
rect 253204 14418 253256 14424
rect 252928 8968 252980 8974
rect 252928 8910 252980 8916
rect 250260 6316 250312 6322
rect 250260 6258 250312 6264
rect 248788 6180 248840 6186
rect 248788 6122 248840 6128
rect 247684 3528 247736 3534
rect 247132 3460 247184 3466
rect 247420 3454 247632 3482
rect 247684 3470 247736 3476
rect 247132 3402 247184 3408
rect 247604 480 247632 3454
rect 248800 480 248828 6122
rect 254136 4962 254164 304234
rect 254228 293282 254256 306206
rect 254216 293276 254268 293282
rect 254216 293218 254268 293224
rect 254124 4956 254176 4962
rect 254124 4898 254176 4904
rect 253480 4140 253532 4146
rect 253480 4082 253532 4088
rect 251180 3528 251232 3534
rect 251180 3470 251232 3476
rect 249984 3460 250036 3466
rect 249984 3402 250036 3408
rect 249996 480 250024 3402
rect 251192 480 251220 3470
rect 252376 3256 252428 3262
rect 252376 3198 252428 3204
rect 252388 480 252416 3198
rect 253492 480 253520 4082
rect 254320 3602 254348 306870
rect 254412 304450 254440 310420
rect 254412 304422 254532 304450
rect 254400 304360 254452 304366
rect 254400 304302 254452 304308
rect 254412 3670 254440 304302
rect 254504 297566 254532 304422
rect 254596 304366 254624 310420
rect 254676 307896 254728 307902
rect 254676 307838 254728 307844
rect 254584 304360 254636 304366
rect 254584 304302 254636 304308
rect 254492 297560 254544 297566
rect 254492 297502 254544 297508
rect 254688 296714 254716 307838
rect 254780 306270 254808 310420
rect 254964 308786 254992 310420
rect 254952 308780 255004 308786
rect 254952 308722 255004 308728
rect 254768 306264 254820 306270
rect 254768 306206 254820 306212
rect 255148 304298 255176 310420
rect 255332 306134 255360 310420
rect 255516 308718 255544 310420
rect 255504 308712 255556 308718
rect 255504 308654 255556 308660
rect 255504 306400 255556 306406
rect 255504 306342 255556 306348
rect 255412 306332 255464 306338
rect 255412 306274 255464 306280
rect 255320 306128 255372 306134
rect 255320 306070 255372 306076
rect 255136 304292 255188 304298
rect 255136 304234 255188 304240
rect 254596 296686 254716 296714
rect 254596 127634 254624 296686
rect 254584 127628 254636 127634
rect 254584 127570 254636 127576
rect 255424 11762 255452 306274
rect 255516 93158 255544 306342
rect 255700 306082 255728 310420
rect 255884 306406 255912 310420
rect 256068 308854 256096 310420
rect 256056 308848 256108 308854
rect 256056 308790 256108 308796
rect 256148 308848 256200 308854
rect 256148 308790 256200 308796
rect 255964 307828 256016 307834
rect 255964 307770 256016 307776
rect 255872 306400 255924 306406
rect 255872 306342 255924 306348
rect 255872 306128 255924 306134
rect 255700 306054 255820 306082
rect 255872 306070 255924 306076
rect 255596 305992 255648 305998
rect 255596 305934 255648 305940
rect 255608 104174 255636 305934
rect 255688 305924 255740 305930
rect 255688 305866 255740 305872
rect 255700 137290 255728 305866
rect 255688 137284 255740 137290
rect 255688 137226 255740 137232
rect 255596 104168 255648 104174
rect 255596 104110 255648 104116
rect 255504 93152 255556 93158
rect 255504 93094 255556 93100
rect 255504 89004 255556 89010
rect 255504 88946 255556 88952
rect 255516 16574 255544 88946
rect 255516 16546 255728 16574
rect 255412 11756 255464 11762
rect 255412 11698 255464 11704
rect 254676 6248 254728 6254
rect 254676 6190 254728 6196
rect 254400 3664 254452 3670
rect 254400 3606 254452 3612
rect 254308 3596 254360 3602
rect 254308 3538 254360 3544
rect 254688 480 254716 6190
rect 255700 3482 255728 16546
rect 255792 6390 255820 306054
rect 255884 291922 255912 306070
rect 255872 291916 255924 291922
rect 255872 291858 255924 291864
rect 255976 13122 256004 307770
rect 256160 305538 256188 308790
rect 256252 305930 256280 310420
rect 256436 306338 256464 310420
rect 256424 306332 256476 306338
rect 256424 306274 256476 306280
rect 256620 305998 256648 310420
rect 256804 306354 256832 310420
rect 256988 307834 257016 310420
rect 257172 308582 257200 310420
rect 257160 308576 257212 308582
rect 257160 308518 257212 308524
rect 256976 307828 257028 307834
rect 256976 307770 257028 307776
rect 256804 306326 257016 306354
rect 256792 306264 256844 306270
rect 256792 306206 256844 306212
rect 256608 305992 256660 305998
rect 256608 305934 256660 305940
rect 256240 305924 256292 305930
rect 256240 305866 256292 305872
rect 256068 305510 256188 305538
rect 256068 156777 256096 305510
rect 256148 303204 256200 303210
rect 256148 303146 256200 303152
rect 256054 156768 256110 156777
rect 256054 156703 256110 156712
rect 256160 152998 256188 303146
rect 256240 303068 256292 303074
rect 256240 303010 256292 303016
rect 256148 152992 256200 152998
rect 256148 152934 256200 152940
rect 256252 152930 256280 303010
rect 256240 152924 256292 152930
rect 256240 152866 256292 152872
rect 256804 91798 256832 306206
rect 256884 306196 256936 306202
rect 256884 306138 256936 306144
rect 256896 95946 256924 306138
rect 256988 306082 257016 306326
rect 257160 306128 257212 306134
rect 256988 306054 257108 306082
rect 257160 306070 257212 306076
rect 256976 305992 257028 305998
rect 256976 305934 257028 305940
rect 256988 138718 257016 305934
rect 257080 140078 257108 306054
rect 257068 140072 257120 140078
rect 257068 140014 257120 140020
rect 256976 138712 257028 138718
rect 256976 138654 257028 138660
rect 256884 95940 256936 95946
rect 256884 95882 256936 95888
rect 256792 91792 256844 91798
rect 256792 91734 256844 91740
rect 257172 26926 257200 306070
rect 257356 305998 257384 310420
rect 257436 308712 257488 308718
rect 257436 308654 257488 308660
rect 257344 305992 257396 305998
rect 257344 305934 257396 305940
rect 257344 305584 257396 305590
rect 257344 305526 257396 305532
rect 257160 26920 257212 26926
rect 257160 26862 257212 26868
rect 256700 14476 256752 14482
rect 256700 14418 256752 14424
rect 255964 13116 256016 13122
rect 255964 13058 256016 13064
rect 255780 6384 255832 6390
rect 255780 6326 255832 6332
rect 255700 3454 255912 3482
rect 255884 480 255912 3454
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 354 256740 14418
rect 257356 6526 257384 305526
rect 257448 155281 257476 308654
rect 257540 306270 257568 310420
rect 257528 306264 257580 306270
rect 257528 306206 257580 306212
rect 257724 306134 257752 310420
rect 257802 308544 257858 308553
rect 257802 308479 257858 308488
rect 257712 306128 257764 306134
rect 257712 306070 257764 306076
rect 257816 302234 257844 308479
rect 257908 306202 257936 310420
rect 257988 308916 258040 308922
rect 257988 308858 258040 308864
rect 257896 306196 257948 306202
rect 257896 306138 257948 306144
rect 258000 305590 258028 308858
rect 258092 306626 258120 310420
rect 258276 309058 258304 310420
rect 258264 309052 258316 309058
rect 258264 308994 258316 309000
rect 258460 307902 258488 310420
rect 258644 308106 258672 310420
rect 258632 308100 258684 308106
rect 258632 308042 258684 308048
rect 258448 307896 258500 307902
rect 258448 307838 258500 307844
rect 258092 306598 258396 306626
rect 258828 306610 258856 310420
rect 258264 306400 258316 306406
rect 258264 306342 258316 306348
rect 258172 306264 258224 306270
rect 258172 306206 258224 306212
rect 257988 305584 258040 305590
rect 257988 305526 258040 305532
rect 257540 302206 257844 302234
rect 257540 158982 257568 302206
rect 257528 158976 257580 158982
rect 257528 158918 257580 158924
rect 257434 155272 257490 155281
rect 257434 155207 257490 155216
rect 258184 105602 258212 306206
rect 258276 130422 258304 306342
rect 258368 141438 258396 306598
rect 258816 306604 258868 306610
rect 258816 306546 258868 306552
rect 259012 306490 259040 310420
rect 258460 306462 259040 306490
rect 258460 149734 258488 306462
rect 259196 306354 259224 310420
rect 258552 306326 259224 306354
rect 258448 149728 258500 149734
rect 258448 149670 258500 149676
rect 258356 141432 258408 141438
rect 258356 141374 258408 141380
rect 258264 130416 258316 130422
rect 258264 130358 258316 130364
rect 258172 105596 258224 105602
rect 258172 105538 258224 105544
rect 258552 90370 258580 306326
rect 259380 306270 259408 310420
rect 259564 306626 259592 310420
rect 259564 306598 259684 306626
rect 259552 306468 259604 306474
rect 259552 306410 259604 306416
rect 259460 306400 259512 306406
rect 259460 306342 259512 306348
rect 259368 306264 259420 306270
rect 259368 306206 259420 306212
rect 258908 303408 258960 303414
rect 258908 303350 258960 303356
rect 258816 303340 258868 303346
rect 258816 303282 258868 303288
rect 258724 303272 258776 303278
rect 258724 303214 258776 303220
rect 258736 153066 258764 303214
rect 258828 153134 258856 303282
rect 258920 153202 258948 303350
rect 258908 153196 258960 153202
rect 258908 153138 258960 153144
rect 258816 153128 258868 153134
rect 258816 153070 258868 153076
rect 258724 153060 258776 153066
rect 258724 153002 258776 153008
rect 259472 108322 259500 306342
rect 259564 116618 259592 306410
rect 259656 306270 259684 306598
rect 259644 306264 259696 306270
rect 259644 306206 259696 306212
rect 259644 306128 259696 306134
rect 259644 306070 259696 306076
rect 259656 129062 259684 306070
rect 259748 141506 259776 310420
rect 259932 306474 259960 310420
rect 259920 306468 259972 306474
rect 259920 306410 259972 306416
rect 260116 306354 260144 310420
rect 260196 307828 260248 307834
rect 260196 307770 260248 307776
rect 259828 306332 259880 306338
rect 259828 306274 259880 306280
rect 259932 306326 260144 306354
rect 259840 144226 259868 306274
rect 259932 148374 259960 306326
rect 260012 306264 260064 306270
rect 260012 306206 260064 306212
rect 260024 174690 260052 306206
rect 260208 296714 260236 307770
rect 260300 306134 260328 310420
rect 260484 306406 260512 310420
rect 260472 306400 260524 306406
rect 260472 306342 260524 306348
rect 260668 306338 260696 310420
rect 260656 306332 260708 306338
rect 260656 306274 260708 306280
rect 260852 306270 260880 310420
rect 260932 306332 260984 306338
rect 260932 306274 260984 306280
rect 260840 306264 260892 306270
rect 260840 306206 260892 306212
rect 260288 306128 260340 306134
rect 260288 306070 260340 306076
rect 260840 306128 260892 306134
rect 260840 306070 260892 306076
rect 260116 296686 260236 296714
rect 260012 174684 260064 174690
rect 260012 174626 260064 174632
rect 259920 148368 259972 148374
rect 259920 148310 259972 148316
rect 259828 144220 259880 144226
rect 259828 144162 259880 144168
rect 260116 142866 260144 296686
rect 260196 144220 260248 144226
rect 260196 144162 260248 144168
rect 260104 142860 260156 142866
rect 260104 142802 260156 142808
rect 259736 141500 259788 141506
rect 259736 141442 259788 141448
rect 259644 129056 259696 129062
rect 259644 128998 259696 129004
rect 259552 116612 259604 116618
rect 259552 116554 259604 116560
rect 259460 108316 259512 108322
rect 259460 108258 259512 108264
rect 260104 108316 260156 108322
rect 260104 108258 260156 108264
rect 258540 90364 258592 90370
rect 258540 90306 258592 90312
rect 259460 15904 259512 15910
rect 259460 15846 259512 15852
rect 257344 6520 257396 6526
rect 257344 6462 257396 6468
rect 258262 3360 258318 3369
rect 258262 3295 258318 3304
rect 258276 480 258304 3295
rect 259472 480 259500 15846
rect 260116 3262 260144 108258
rect 260208 4146 260236 144162
rect 260852 19990 260880 306070
rect 260944 101454 260972 306274
rect 261036 102814 261064 310420
rect 261220 306513 261248 310420
rect 261404 306626 261432 310420
rect 261312 306598 261432 306626
rect 261206 306504 261262 306513
rect 261206 306439 261262 306448
rect 261116 306400 261168 306406
rect 261312 306354 261340 306598
rect 261116 306342 261168 306348
rect 261128 122126 261156 306342
rect 261220 306326 261340 306354
rect 261588 306338 261616 310420
rect 261576 306332 261628 306338
rect 261220 123486 261248 306326
rect 261576 306274 261628 306280
rect 261300 306264 261352 306270
rect 261772 306218 261800 310420
rect 261956 306406 261984 310420
rect 261944 306400 261996 306406
rect 261944 306342 261996 306348
rect 261300 306206 261352 306212
rect 261312 145586 261340 306206
rect 261404 306190 261800 306218
rect 261404 146946 261432 306190
rect 262140 306134 262168 310420
rect 262324 307834 262352 310420
rect 262312 307828 262364 307834
rect 262312 307770 262364 307776
rect 262312 306400 262364 306406
rect 262508 306354 262536 310420
rect 262312 306342 262364 306348
rect 262128 306128 262180 306134
rect 261482 306096 261538 306105
rect 262128 306070 262180 306076
rect 261482 306031 261538 306040
rect 261496 152522 261524 306031
rect 261668 303476 261720 303482
rect 261668 303418 261720 303424
rect 261576 302932 261628 302938
rect 261576 302874 261628 302880
rect 261588 155038 261616 302874
rect 261680 157321 261708 303418
rect 261666 157312 261722 157321
rect 261666 157247 261722 157256
rect 261576 155032 261628 155038
rect 261576 154974 261628 154980
rect 261484 152516 261536 152522
rect 261484 152458 261536 152464
rect 261392 146940 261444 146946
rect 261392 146882 261444 146888
rect 261300 145580 261352 145586
rect 261300 145522 261352 145528
rect 261208 123480 261260 123486
rect 261208 123422 261260 123428
rect 261116 122120 261168 122126
rect 261116 122062 261168 122068
rect 262324 120766 262352 306342
rect 262416 306326 262536 306354
rect 262588 306332 262640 306338
rect 262416 134570 262444 306326
rect 262588 306274 262640 306280
rect 262496 306264 262548 306270
rect 262496 306206 262548 306212
rect 262508 145654 262536 306206
rect 262600 151094 262628 306274
rect 262692 156641 262720 310420
rect 262876 306338 262904 310420
rect 263060 306406 263088 310420
rect 263048 306400 263100 306406
rect 263048 306342 263100 306348
rect 262864 306332 262916 306338
rect 262864 306274 262916 306280
rect 263244 296714 263272 310420
rect 263428 306270 263456 310420
rect 263612 308310 263640 310420
rect 263796 308394 263824 310420
rect 263980 308718 264008 310420
rect 263968 308712 264020 308718
rect 263968 308654 264020 308660
rect 264164 308428 264192 310420
rect 263704 308366 263824 308394
rect 263888 308400 264192 308428
rect 263600 308304 263652 308310
rect 263600 308246 263652 308252
rect 263416 306264 263468 306270
rect 263416 306206 263468 306212
rect 262784 296686 263272 296714
rect 262678 156632 262734 156641
rect 262678 156567 262734 156576
rect 262588 151088 262640 151094
rect 262588 151030 262640 151036
rect 262496 145648 262548 145654
rect 262496 145590 262548 145596
rect 262404 134564 262456 134570
rect 262404 134506 262456 134512
rect 262312 120760 262364 120766
rect 262312 120702 262364 120708
rect 261024 102808 261076 102814
rect 261024 102750 261076 102756
rect 260932 101448 260984 101454
rect 260932 101390 260984 101396
rect 262784 100026 262812 296686
rect 262772 100020 262824 100026
rect 262772 99962 262824 99968
rect 263704 98666 263732 308366
rect 263784 308236 263836 308242
rect 263784 308178 263836 308184
rect 263796 117978 263824 308178
rect 263888 119406 263916 308400
rect 263968 308304 264020 308310
rect 263968 308246 264020 308252
rect 263980 133210 264008 308246
rect 264348 307034 264376 310420
rect 264072 307006 264376 307034
rect 264072 135930 264100 307006
rect 264532 306898 264560 310420
rect 264612 308440 264664 308446
rect 264612 308382 264664 308388
rect 264164 306870 264560 306898
rect 264164 149802 264192 306870
rect 264624 306762 264652 308382
rect 264716 308242 264744 310420
rect 264704 308236 264756 308242
rect 264704 308178 264756 308184
rect 264256 306734 264652 306762
rect 264152 149796 264204 149802
rect 264152 149738 264204 149744
rect 264060 135924 264112 135930
rect 264060 135866 264112 135872
rect 263968 133204 264020 133210
rect 263968 133146 264020 133152
rect 263876 119400 263928 119406
rect 263876 119342 263928 119348
rect 263784 117972 263836 117978
rect 263784 117914 263836 117920
rect 263692 98660 263744 98666
rect 263692 98602 263744 98608
rect 260840 19984 260892 19990
rect 260840 19926 260892 19932
rect 261760 6928 261812 6934
rect 261760 6870 261812 6876
rect 260196 4140 260248 4146
rect 260196 4082 260248 4088
rect 260656 3392 260708 3398
rect 260656 3334 260708 3340
rect 260104 3256 260156 3262
rect 260104 3198 260156 3204
rect 260668 480 260696 3334
rect 261772 480 261800 6870
rect 264256 3806 264284 306734
rect 264426 303512 264482 303521
rect 264426 303447 264482 303456
rect 264336 303000 264388 303006
rect 264336 302942 264388 302948
rect 264348 155106 264376 302942
rect 264440 155961 264468 303447
rect 264900 296714 264928 310420
rect 265084 308446 265112 310420
rect 265072 308440 265124 308446
rect 265072 308382 265124 308388
rect 265164 308440 265216 308446
rect 265164 308382 265216 308388
rect 265072 308304 265124 308310
rect 265072 308246 265124 308252
rect 264532 296686 264928 296714
rect 264426 155952 264482 155961
rect 264426 155887 264482 155896
rect 264336 155100 264388 155106
rect 264336 155042 264388 155048
rect 264532 21418 264560 296686
rect 265084 113830 265112 308246
rect 265176 115258 265204 308382
rect 265268 308156 265296 310420
rect 265452 308446 265480 310420
rect 265440 308440 265492 308446
rect 265636 308394 265664 310420
rect 265440 308382 265492 308388
rect 265544 308366 265664 308394
rect 265440 308168 265492 308174
rect 265268 308128 265388 308156
rect 265256 308032 265308 308038
rect 265256 307974 265308 307980
rect 265268 138786 265296 307974
rect 265360 140146 265388 308128
rect 265440 308110 265492 308116
rect 265452 153882 265480 308110
rect 265440 153876 265492 153882
rect 265440 153818 265492 153824
rect 265348 140140 265400 140146
rect 265348 140082 265400 140088
rect 265256 138780 265308 138786
rect 265256 138722 265308 138728
rect 265164 115252 265216 115258
rect 265164 115194 265216 115200
rect 265072 113824 265124 113830
rect 265072 113766 265124 113772
rect 264520 21412 264572 21418
rect 264520 21354 264572 21360
rect 265544 5030 265572 308366
rect 265820 308038 265848 310420
rect 266004 308310 266032 310420
rect 265992 308304 266044 308310
rect 265992 308246 266044 308252
rect 266188 308174 266216 310420
rect 266372 308310 266400 310420
rect 266452 309052 266504 309058
rect 266452 308994 266504 309000
rect 266464 308922 266492 308994
rect 266452 308916 266504 308922
rect 266452 308858 266504 308864
rect 266452 308440 266504 308446
rect 266452 308382 266504 308388
rect 266360 308304 266412 308310
rect 266360 308246 266412 308252
rect 266176 308168 266228 308174
rect 266176 308110 266228 308116
rect 265808 308032 265860 308038
rect 265808 307974 265860 307980
rect 265624 307828 265676 307834
rect 265624 307770 265676 307776
rect 265636 131850 265664 307770
rect 265714 303376 265770 303385
rect 265714 303311 265770 303320
rect 265728 155378 265756 303311
rect 265716 155372 265768 155378
rect 265716 155314 265768 155320
rect 265624 131844 265676 131850
rect 265624 131786 265676 131792
rect 266464 6458 266492 308382
rect 266556 308292 266584 310420
rect 266740 308394 266768 310420
rect 266924 308446 266952 310420
rect 267108 309074 267136 310420
rect 267016 309046 267136 309074
rect 266912 308440 266964 308446
rect 266740 308366 266860 308394
rect 266912 308382 266964 308388
rect 266556 308264 266768 308292
rect 266636 308168 266688 308174
rect 266636 308110 266688 308116
rect 266544 308100 266596 308106
rect 266544 308042 266596 308048
rect 266556 7682 266584 308042
rect 266648 112470 266676 308110
rect 266740 124914 266768 308264
rect 266832 173194 266860 308366
rect 266912 308304 266964 308310
rect 266912 308246 266964 308252
rect 266820 173188 266872 173194
rect 266820 173130 266872 173136
rect 266728 124908 266780 124914
rect 266728 124850 266780 124856
rect 266636 112464 266688 112470
rect 266636 112406 266688 112412
rect 266544 7676 266596 7682
rect 266544 7618 266596 7624
rect 266452 6452 266504 6458
rect 266452 6394 266504 6400
rect 266924 5098 266952 308246
rect 267016 308174 267044 309046
rect 267096 308916 267148 308922
rect 267096 308858 267148 308864
rect 267004 308168 267056 308174
rect 267004 308110 267056 308116
rect 267004 305652 267056 305658
rect 267004 305594 267056 305600
rect 267016 155242 267044 305594
rect 267108 159186 267136 308858
rect 267292 308854 267320 310420
rect 267476 309058 267504 310420
rect 267464 309052 267516 309058
rect 267464 308994 267516 309000
rect 267280 308848 267332 308854
rect 267280 308790 267332 308796
rect 267660 308106 267688 310420
rect 267844 308666 267872 310420
rect 267844 308638 267964 308666
rect 267832 308508 267884 308514
rect 267832 308450 267884 308456
rect 267740 308440 267792 308446
rect 267740 308382 267792 308388
rect 267648 308100 267700 308106
rect 267648 308042 267700 308048
rect 267188 303136 267240 303142
rect 267188 303078 267240 303084
rect 267096 159180 267148 159186
rect 267096 159122 267148 159128
rect 267004 155236 267056 155242
rect 267004 155178 267056 155184
rect 267200 155174 267228 303078
rect 267188 155168 267240 155174
rect 267188 155110 267240 155116
rect 267004 134564 267056 134570
rect 267004 134506 267056 134512
rect 266912 5092 266964 5098
rect 266912 5034 266964 5040
rect 265532 5024 265584 5030
rect 265532 4966 265584 4972
rect 265348 4956 265400 4962
rect 265348 4898 265400 4904
rect 264244 3800 264296 3806
rect 264244 3742 264296 3748
rect 264152 3664 264204 3670
rect 264152 3606 264204 3612
rect 262956 3596 263008 3602
rect 262956 3538 263008 3544
rect 262968 480 262996 3538
rect 264164 480 264192 3606
rect 265360 480 265388 4898
rect 266544 3936 266596 3942
rect 266544 3878 266596 3884
rect 266556 480 266584 3878
rect 267016 3602 267044 134506
rect 267752 111110 267780 308382
rect 267844 126274 267872 308450
rect 267936 308310 267964 308638
rect 267924 308304 267976 308310
rect 267924 308246 267976 308252
rect 267924 308168 267976 308174
rect 267924 308110 267976 308116
rect 267936 133278 267964 308110
rect 268028 134638 268056 310420
rect 268212 308514 268240 310420
rect 268200 308508 268252 308514
rect 268200 308450 268252 308456
rect 268396 308394 268424 310420
rect 268212 308366 268424 308394
rect 268108 306604 268160 306610
rect 268108 306546 268160 306552
rect 268120 149870 268148 306546
rect 268212 151162 268240 308366
rect 268292 308304 268344 308310
rect 268292 308246 268344 308252
rect 268304 155417 268332 308246
rect 268384 308236 268436 308242
rect 268384 308178 268436 308184
rect 268290 155408 268346 155417
rect 268290 155343 268346 155352
rect 268200 151156 268252 151162
rect 268200 151098 268252 151104
rect 268108 149864 268160 149870
rect 268108 149806 268160 149812
rect 268016 134632 268068 134638
rect 268016 134574 268068 134580
rect 267924 133272 267976 133278
rect 267924 133214 267976 133220
rect 267832 126268 267884 126274
rect 267832 126210 267884 126216
rect 267740 111104 267792 111110
rect 267740 111046 267792 111052
rect 267740 17332 267792 17338
rect 267740 17274 267792 17280
rect 267004 3596 267056 3602
rect 267004 3538 267056 3544
rect 267096 3596 267148 3602
rect 267096 3538 267148 3544
rect 267108 3398 267136 3538
rect 267096 3392 267148 3398
rect 267096 3334 267148 3340
rect 267752 480 267780 17274
rect 268396 5302 268424 308178
rect 268580 308174 268608 310420
rect 268764 308446 268792 310420
rect 268752 308440 268804 308446
rect 268752 308382 268804 308388
rect 268568 308168 268620 308174
rect 268568 308110 268620 308116
rect 268948 306610 268976 310420
rect 269132 308310 269160 310420
rect 269316 308530 269344 310420
rect 269500 308530 269528 310420
rect 269224 308502 269344 308530
rect 269408 308502 269528 308530
rect 269120 308304 269172 308310
rect 269120 308246 269172 308252
rect 269224 307834 269252 308502
rect 269304 308440 269356 308446
rect 269304 308382 269356 308388
rect 269212 307828 269264 307834
rect 269212 307770 269264 307776
rect 269212 307692 269264 307698
rect 269212 307634 269264 307640
rect 268936 306604 268988 306610
rect 268936 306546 268988 306552
rect 268474 151056 268530 151065
rect 268474 150991 268530 151000
rect 268384 5296 268436 5302
rect 268384 5238 268436 5244
rect 268488 3466 268516 150991
rect 268568 133204 268620 133210
rect 268568 133146 268620 133152
rect 268580 3534 268608 133146
rect 269224 17270 269252 307634
rect 269316 109750 269344 308382
rect 269408 308174 269436 308502
rect 269684 308394 269712 310420
rect 269868 308446 269896 310420
rect 269500 308366 269712 308394
rect 269856 308440 269908 308446
rect 269856 308382 269908 308388
rect 269396 308168 269448 308174
rect 269396 308110 269448 308116
rect 269396 308032 269448 308038
rect 269396 307974 269448 307980
rect 269408 130490 269436 307974
rect 269500 131782 269528 308366
rect 269580 308304 269632 308310
rect 270052 308258 270080 310420
rect 269580 308246 269632 308252
rect 269592 144294 269620 308246
rect 269684 308230 270080 308258
rect 269684 153950 269712 308230
rect 269948 308168 270000 308174
rect 269948 308110 270000 308116
rect 269764 307828 269816 307834
rect 269764 307770 269816 307776
rect 269672 153944 269724 153950
rect 269672 153886 269724 153892
rect 269580 144288 269632 144294
rect 269580 144230 269632 144236
rect 269488 131776 269540 131782
rect 269488 131718 269540 131724
rect 269396 130484 269448 130490
rect 269396 130426 269448 130432
rect 269304 109744 269356 109750
rect 269304 109686 269356 109692
rect 269212 17264 269264 17270
rect 269212 17206 269264 17212
rect 269776 6934 269804 307770
rect 269856 305788 269908 305794
rect 269856 305730 269908 305736
rect 269868 158409 269896 305730
rect 269854 158400 269910 158409
rect 269854 158335 269910 158344
rect 269856 111104 269908 111110
rect 269856 111046 269908 111052
rect 269764 6928 269816 6934
rect 269764 6870 269816 6876
rect 269868 3942 269896 111046
rect 269960 5166 269988 308110
rect 270236 308038 270264 310420
rect 270224 308032 270276 308038
rect 270224 307974 270276 307980
rect 270420 307698 270448 310420
rect 270500 308508 270552 308514
rect 270500 308450 270552 308456
rect 270408 307692 270460 307698
rect 270408 307634 270460 307640
rect 270040 305720 270092 305726
rect 270040 305662 270092 305668
rect 270052 158273 270080 305662
rect 270038 158264 270094 158273
rect 270038 158199 270094 158208
rect 270512 106962 270540 308450
rect 270604 308281 270632 310420
rect 270684 308372 270736 308378
rect 270684 308314 270736 308320
rect 270590 308272 270646 308281
rect 270590 308207 270646 308216
rect 270592 307420 270644 307426
rect 270592 307362 270644 307368
rect 270604 129130 270632 307362
rect 270696 141574 270724 308314
rect 270788 142934 270816 310420
rect 270972 307426 271000 310420
rect 270960 307420 271012 307426
rect 270960 307362 271012 307368
rect 271156 306898 271184 310420
rect 271236 308440 271288 308446
rect 271236 308382 271288 308388
rect 270880 306870 271184 306898
rect 270880 147014 270908 306870
rect 270960 306808 271012 306814
rect 270960 306750 271012 306756
rect 270972 156913 271000 306750
rect 271248 296714 271276 308382
rect 271340 308378 271368 310420
rect 271524 308514 271552 310420
rect 271512 308508 271564 308514
rect 271512 308450 271564 308456
rect 271328 308372 271380 308378
rect 271328 308314 271380 308320
rect 271708 306814 271736 310420
rect 271892 308446 271920 310420
rect 271880 308440 271932 308446
rect 271880 308382 271932 308388
rect 271972 308372 272024 308378
rect 271972 308314 272024 308320
rect 271696 306808 271748 306814
rect 271696 306750 271748 306756
rect 271788 306264 271840 306270
rect 271788 306206 271840 306212
rect 271696 306128 271748 306134
rect 271696 306070 271748 306076
rect 271604 303544 271656 303550
rect 271604 303486 271656 303492
rect 271156 296686 271276 296714
rect 270958 156904 271014 156913
rect 270958 156839 271014 156848
rect 270868 147008 270920 147014
rect 270868 146950 270920 146956
rect 270960 146940 271012 146946
rect 270960 146882 271012 146888
rect 270776 142928 270828 142934
rect 270776 142870 270828 142876
rect 270684 141568 270736 141574
rect 270684 141510 270736 141516
rect 270592 129124 270644 129130
rect 270592 129066 270644 129072
rect 270500 106956 270552 106962
rect 270500 106898 270552 106904
rect 269948 5160 270000 5166
rect 269948 5102 270000 5108
rect 269856 3936 269908 3942
rect 269856 3878 269908 3884
rect 268568 3528 268620 3534
rect 268568 3470 268620 3476
rect 268844 3528 268896 3534
rect 268844 3470 268896 3476
rect 268476 3460 268528 3466
rect 268476 3402 268528 3408
rect 268856 480 268884 3470
rect 270040 3460 270092 3466
rect 270040 3402 270092 3408
rect 270052 480 270080 3402
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270972 354 271000 146882
rect 271156 127702 271184 296686
rect 271616 158409 271644 303486
rect 271602 158400 271658 158409
rect 271602 158335 271658 158344
rect 271616 158030 271644 158335
rect 271708 158273 271736 306070
rect 271694 158264 271750 158273
rect 271694 158199 271750 158208
rect 271708 158098 271736 158199
rect 271696 158092 271748 158098
rect 271696 158034 271748 158040
rect 271604 158024 271656 158030
rect 271604 157966 271656 157972
rect 271328 157888 271380 157894
rect 271328 157830 271380 157836
rect 271420 157888 271472 157894
rect 271420 157830 271472 157836
rect 271340 157554 271368 157830
rect 271432 157729 271460 157830
rect 271418 157720 271474 157729
rect 271418 157655 271474 157664
rect 271328 157548 271380 157554
rect 271328 157490 271380 157496
rect 271800 154562 271828 306206
rect 271788 154556 271840 154562
rect 271788 154498 271840 154504
rect 271800 154154 271828 154498
rect 271788 154148 271840 154154
rect 271788 154090 271840 154096
rect 271236 152516 271288 152522
rect 271236 152458 271288 152464
rect 271144 127696 271196 127702
rect 271144 127638 271196 127644
rect 271248 3602 271276 152458
rect 271984 18630 272012 308314
rect 272076 130558 272104 310420
rect 272156 308440 272208 308446
rect 272156 308382 272208 308388
rect 272168 140214 272196 308382
rect 272260 308310 272288 310420
rect 272444 308394 272472 310420
rect 272352 308366 272472 308394
rect 272248 308304 272300 308310
rect 272248 308246 272300 308252
rect 272248 308168 272300 308174
rect 272248 308110 272300 308116
rect 272260 143002 272288 308110
rect 272352 154018 272380 308366
rect 272432 308304 272484 308310
rect 272432 308246 272484 308252
rect 272340 154012 272392 154018
rect 272340 153954 272392 153960
rect 272248 142996 272300 143002
rect 272248 142938 272300 142944
rect 272156 140208 272208 140214
rect 272156 140150 272208 140156
rect 272064 130552 272116 130558
rect 272064 130494 272116 130500
rect 271972 18624 272024 18630
rect 271972 18566 272024 18572
rect 272444 5234 272472 308246
rect 272628 308174 272656 310420
rect 272812 308242 272840 310420
rect 272996 308446 273024 310420
rect 272984 308440 273036 308446
rect 272984 308382 273036 308388
rect 273180 308378 273208 310420
rect 273168 308372 273220 308378
rect 273168 308314 273220 308320
rect 272800 308236 272852 308242
rect 272800 308178 272852 308184
rect 272616 308168 272668 308174
rect 272616 308110 272668 308116
rect 273364 307873 273392 310420
rect 273548 308009 273576 310420
rect 273534 308000 273590 308009
rect 273534 307935 273590 307944
rect 273350 307864 273406 307873
rect 273350 307799 273406 307808
rect 273260 306400 273312 306406
rect 273732 306354 273760 310420
rect 273260 306342 273312 306348
rect 272616 305924 272668 305930
rect 272616 305866 272668 305872
rect 272524 305856 272576 305862
rect 272524 305798 272576 305804
rect 272536 156534 272564 305798
rect 272524 156528 272576 156534
rect 272524 156470 272576 156476
rect 272628 156466 272656 305866
rect 273168 246696 273220 246702
rect 273168 246638 273220 246644
rect 272616 156460 272668 156466
rect 272616 156402 272668 156408
rect 273180 154562 273208 246638
rect 272708 154556 272760 154562
rect 272708 154498 272760 154504
rect 273168 154556 273220 154562
rect 273168 154498 273220 154504
rect 272720 153814 272748 154498
rect 272708 153808 272760 153814
rect 272708 153750 272760 153756
rect 273272 105670 273300 306342
rect 273352 306332 273404 306338
rect 273352 306274 273404 306280
rect 273456 306326 273760 306354
rect 273364 126342 273392 306274
rect 273456 144362 273484 306326
rect 273916 306218 273944 310420
rect 273996 307828 274048 307834
rect 273996 307770 274048 307776
rect 273548 306190 273944 306218
rect 273548 145722 273576 306190
rect 273628 306060 273680 306066
rect 273628 306002 273680 306008
rect 273640 155553 273668 306002
rect 274008 302234 274036 307770
rect 274100 306338 274128 310420
rect 274284 306406 274312 310420
rect 274272 306400 274324 306406
rect 274272 306342 274324 306348
rect 274088 306332 274140 306338
rect 274088 306274 274140 306280
rect 274468 306066 274496 310420
rect 274548 308644 274600 308650
rect 274548 308586 274600 308592
rect 274456 306060 274508 306066
rect 274456 306002 274508 306008
rect 274560 305674 274588 308586
rect 274652 307873 274680 310420
rect 274836 308009 274864 310420
rect 274822 308000 274878 308009
rect 274822 307935 274878 307944
rect 274638 307864 274694 307873
rect 275020 307834 275048 310420
rect 274638 307799 274694 307808
rect 275008 307828 275060 307834
rect 275008 307770 275060 307776
rect 274732 306400 274784 306406
rect 275204 306354 275232 310420
rect 274732 306342 274784 306348
rect 274560 305646 274680 305674
rect 274548 305516 274600 305522
rect 274548 305458 274600 305464
rect 274364 305448 274416 305454
rect 274364 305390 274416 305396
rect 273916 302206 274036 302234
rect 273720 157276 273772 157282
rect 273720 157218 273772 157224
rect 273732 156806 273760 157218
rect 273720 156800 273772 156806
rect 273720 156742 273772 156748
rect 273626 155544 273682 155553
rect 273626 155479 273682 155488
rect 273916 148442 273944 302206
rect 274272 246764 274324 246770
rect 274272 246706 274324 246712
rect 274284 161474 274312 246706
rect 274192 161446 274312 161474
rect 274192 157282 274220 161446
rect 274376 158234 274404 305390
rect 274560 303634 274588 305458
rect 274468 303606 274588 303634
rect 274364 158228 274416 158234
rect 274364 158170 274416 158176
rect 274376 157865 274404 158170
rect 274468 158166 274496 303606
rect 274652 303498 274680 305646
rect 274560 303470 274680 303498
rect 274456 158160 274508 158166
rect 274454 158128 274456 158137
rect 274508 158128 274510 158137
rect 274454 158063 274510 158072
rect 274362 157856 274418 157865
rect 274362 157791 274418 157800
rect 274180 157276 274232 157282
rect 274180 157218 274232 157224
rect 274560 156874 274588 303470
rect 274638 157584 274694 157593
rect 274638 157519 274640 157528
rect 274692 157519 274694 157528
rect 274640 157490 274692 157496
rect 274548 156868 274600 156874
rect 274548 156810 274600 156816
rect 274640 155780 274692 155786
rect 274640 155722 274692 155728
rect 274652 155310 274680 155722
rect 274640 155304 274692 155310
rect 274640 155246 274692 155252
rect 273904 148436 273956 148442
rect 273904 148378 273956 148384
rect 273996 148368 274048 148374
rect 273996 148310 274048 148316
rect 273536 145716 273588 145722
rect 273536 145658 273588 145664
rect 273904 145580 273956 145586
rect 273904 145522 273956 145528
rect 273444 144356 273496 144362
rect 273444 144298 273496 144304
rect 273352 126336 273404 126342
rect 273352 126278 273404 126284
rect 273260 105664 273312 105670
rect 273260 105606 273312 105612
rect 272432 5228 272484 5234
rect 272432 5170 272484 5176
rect 273916 3670 273944 145522
rect 273904 3664 273956 3670
rect 273904 3606 273956 3612
rect 271236 3596 271288 3602
rect 271236 3538 271288 3544
rect 274008 3466 274036 148310
rect 274088 138712 274140 138718
rect 274088 138654 274140 138660
rect 274100 3534 274128 138654
rect 274744 104242 274772 306342
rect 274824 306332 274876 306338
rect 274824 306274 274876 306280
rect 274928 306326 275232 306354
rect 274836 124982 274864 306274
rect 274928 137358 274956 306326
rect 275388 306218 275416 310420
rect 275468 307828 275520 307834
rect 275468 307770 275520 307776
rect 275008 306196 275060 306202
rect 275008 306138 275060 306144
rect 275112 306190 275416 306218
rect 275020 154086 275048 306138
rect 275008 154080 275060 154086
rect 275008 154022 275060 154028
rect 274916 137352 274968 137358
rect 274916 137294 274968 137300
rect 274824 124976 274876 124982
rect 274824 124918 274876 124924
rect 274732 104236 274784 104242
rect 274732 104178 274784 104184
rect 275112 10402 275140 306190
rect 275284 305992 275336 305998
rect 275284 305934 275336 305940
rect 275296 156602 275324 305934
rect 275376 305584 275428 305590
rect 275376 305526 275428 305532
rect 275388 156670 275416 305526
rect 275480 159497 275508 307770
rect 275572 306202 275600 310420
rect 275756 306338 275784 310420
rect 275940 306406 275968 310420
rect 276124 307834 276152 310420
rect 276112 307828 276164 307834
rect 276112 307770 276164 307776
rect 275928 306400 275980 306406
rect 275928 306342 275980 306348
rect 276204 306400 276256 306406
rect 276204 306342 276256 306348
rect 276308 306354 276336 310420
rect 276492 306354 276520 310420
rect 275744 306332 275796 306338
rect 275744 306274 275796 306280
rect 276112 306332 276164 306338
rect 276112 306274 276164 306280
rect 275560 306196 275612 306202
rect 275560 306138 275612 306144
rect 275928 250844 275980 250850
rect 275928 250786 275980 250792
rect 275836 246832 275888 246838
rect 275836 246774 275888 246780
rect 275466 159488 275522 159497
rect 275466 159423 275522 159432
rect 275376 156664 275428 156670
rect 275376 156606 275428 156612
rect 275284 156596 275336 156602
rect 275284 156538 275336 156544
rect 275848 155786 275876 246774
rect 275940 157593 275968 250786
rect 276018 158536 276074 158545
rect 276018 158471 276074 158480
rect 276032 157962 276060 158471
rect 276020 157956 276072 157962
rect 276020 157898 276072 157904
rect 275926 157584 275982 157593
rect 275926 157519 275982 157528
rect 275836 155780 275888 155786
rect 275836 155722 275888 155728
rect 275284 124908 275336 124914
rect 275284 124850 275336 124856
rect 275100 10396 275152 10402
rect 275100 10338 275152 10344
rect 274824 10328 274876 10334
rect 274824 10270 274876 10276
rect 274088 3528 274140 3534
rect 274088 3470 274140 3476
rect 273996 3460 274048 3466
rect 273996 3402 274048 3408
rect 272432 3256 272484 3262
rect 272432 3198 272484 3204
rect 272444 480 272472 3198
rect 273628 2848 273680 2854
rect 273628 2790 273680 2796
rect 273640 480 273668 2790
rect 274836 480 274864 10270
rect 275296 3262 275324 124850
rect 276124 6594 276152 306274
rect 276216 89214 276244 306342
rect 276308 306326 276428 306354
rect 276492 306326 276612 306354
rect 276676 306338 276704 310420
rect 276296 306060 276348 306066
rect 276296 306002 276348 306008
rect 276204 89208 276256 89214
rect 276204 89150 276256 89156
rect 276308 89146 276336 306002
rect 276296 89140 276348 89146
rect 276296 89082 276348 89088
rect 276400 89078 276428 306326
rect 276480 306196 276532 306202
rect 276480 306138 276532 306144
rect 276492 174554 276520 306138
rect 276480 174548 276532 174554
rect 276480 174490 276532 174496
rect 276388 89072 276440 89078
rect 276388 89014 276440 89020
rect 276584 6662 276612 306326
rect 276664 306332 276716 306338
rect 276664 306274 276716 306280
rect 276860 306066 276888 310420
rect 277044 306202 277072 310420
rect 277124 308576 277176 308582
rect 277124 308518 277176 308524
rect 277032 306196 277084 306202
rect 277032 306138 277084 306144
rect 276848 306060 276900 306066
rect 276848 306002 276900 306008
rect 277136 302234 277164 308518
rect 277228 306406 277256 310420
rect 277308 308508 277360 308514
rect 277308 308450 277360 308456
rect 277216 306400 277268 306406
rect 277216 306342 277268 306348
rect 277136 302206 277256 302234
rect 277124 300348 277176 300354
rect 277124 300290 277176 300296
rect 277032 246968 277084 246974
rect 277032 246910 277084 246916
rect 277044 158545 277072 246910
rect 277030 158536 277086 158545
rect 277030 158471 277086 158480
rect 277136 156942 277164 300290
rect 277228 157010 277256 302206
rect 277216 157004 277268 157010
rect 277216 156946 277268 156952
rect 277124 156936 277176 156942
rect 277124 156878 277176 156884
rect 277320 155446 277348 308450
rect 277412 307873 277440 310420
rect 277398 307864 277454 307873
rect 277398 307799 277454 307808
rect 277596 306542 277624 310420
rect 277780 307018 277808 310420
rect 277768 307012 277820 307018
rect 277768 306954 277820 306960
rect 277676 306808 277728 306814
rect 277676 306750 277728 306756
rect 277584 306536 277636 306542
rect 277584 306478 277636 306484
rect 277492 306468 277544 306474
rect 277492 306410 277544 306416
rect 277308 155440 277360 155446
rect 277308 155382 277360 155388
rect 276572 6656 276624 6662
rect 276572 6598 276624 6604
rect 276112 6588 276164 6594
rect 276112 6530 276164 6536
rect 277504 4894 277532 306410
rect 277584 306332 277636 306338
rect 277584 306274 277636 306280
rect 277596 6186 277624 306274
rect 277688 6730 277716 306750
rect 277860 306536 277912 306542
rect 277860 306478 277912 306484
rect 277768 306060 277820 306066
rect 277768 306002 277820 306008
rect 277780 22778 277808 306002
rect 277872 89282 277900 306478
rect 277964 306218 277992 310420
rect 278148 306474 278176 310420
rect 278228 307896 278280 307902
rect 278228 307838 278280 307844
rect 278136 306468 278188 306474
rect 278136 306410 278188 306416
rect 277964 306190 278176 306218
rect 278044 305380 278096 305386
rect 278044 305322 278096 305328
rect 277952 305312 278004 305318
rect 277952 305254 278004 305260
rect 277964 174622 277992 305254
rect 277952 174616 278004 174622
rect 277952 174558 278004 174564
rect 277950 158672 278006 158681
rect 277950 158607 278006 158616
rect 277964 157894 277992 158607
rect 277952 157888 278004 157894
rect 277952 157830 278004 157836
rect 277860 89276 277912 89282
rect 277860 89218 277912 89224
rect 278056 89010 278084 305322
rect 278044 89004 278096 89010
rect 278044 88946 278096 88952
rect 277768 22772 277820 22778
rect 277768 22714 277820 22720
rect 278044 11620 278096 11626
rect 278044 11562 278096 11568
rect 277676 6724 277728 6730
rect 277676 6666 277728 6672
rect 277584 6180 277636 6186
rect 277584 6122 277636 6128
rect 277492 4888 277544 4894
rect 277492 4830 277544 4836
rect 277124 3528 277176 3534
rect 277124 3470 277176 3476
rect 278056 3482 278084 11562
rect 278148 3738 278176 306190
rect 278240 305386 278268 307838
rect 278228 305380 278280 305386
rect 278228 305322 278280 305328
rect 278332 305318 278360 310420
rect 278516 306066 278544 310420
rect 278700 306338 278728 310420
rect 278884 307873 278912 310420
rect 278870 307864 278926 307873
rect 278870 307799 278926 307808
rect 278964 306468 279016 306474
rect 278964 306410 279016 306416
rect 278688 306332 278740 306338
rect 278688 306274 278740 306280
rect 278504 306060 278556 306066
rect 278504 306002 278556 306008
rect 278596 306060 278648 306066
rect 278596 306002 278648 306008
rect 278608 305590 278636 306002
rect 278596 305584 278648 305590
rect 278596 305526 278648 305532
rect 278320 305312 278372 305318
rect 278320 305254 278372 305260
rect 278872 304700 278924 304706
rect 278872 304642 278924 304648
rect 278596 248192 278648 248198
rect 278596 248134 278648 248140
rect 278608 155582 278636 248134
rect 278688 248124 278740 248130
rect 278688 248066 278740 248072
rect 278596 155576 278648 155582
rect 278596 155518 278648 155524
rect 278700 154222 278728 248066
rect 278688 154216 278740 154222
rect 278688 154158 278740 154164
rect 278884 14482 278912 304642
rect 278976 108322 279004 306410
rect 279068 133210 279096 310420
rect 279252 306474 279280 310420
rect 279240 306468 279292 306474
rect 279240 306410 279292 306416
rect 279436 306354 279464 310420
rect 279160 306326 279464 306354
rect 279160 144226 279188 306326
rect 279620 306082 279648 310420
rect 279804 307902 279832 310420
rect 279792 307896 279844 307902
rect 279792 307838 279844 307844
rect 279884 307896 279936 307902
rect 279884 307838 279936 307844
rect 279700 307828 279752 307834
rect 279700 307770 279752 307776
rect 279252 306054 279648 306082
rect 279148 144220 279200 144226
rect 279148 144162 279200 144168
rect 279056 133204 279108 133210
rect 279056 133146 279108 133152
rect 278964 108316 279016 108322
rect 278964 108258 279016 108264
rect 278964 88800 279016 88806
rect 278964 88742 279016 88748
rect 278976 16574 279004 88742
rect 278976 16546 279096 16574
rect 278872 14476 278924 14482
rect 278872 14418 278924 14424
rect 278688 4412 278740 4418
rect 278688 4354 278740 4360
rect 278136 3732 278188 3738
rect 278136 3674 278188 3680
rect 276020 3460 276072 3466
rect 276020 3402 276072 3408
rect 275284 3256 275336 3262
rect 275284 3198 275336 3204
rect 276032 480 276060 3402
rect 277136 480 277164 3470
rect 278056 3454 278360 3482
rect 278332 480 278360 3454
rect 278700 2854 278728 4354
rect 278688 2848 278740 2854
rect 278688 2790 278740 2796
rect 271206 354 271318 480
rect 270972 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 279252 6254 279280 306054
rect 279424 305584 279476 305590
rect 279424 305526 279476 305532
rect 279240 6248 279292 6254
rect 279240 6190 279292 6196
rect 279436 4962 279464 305526
rect 279712 302234 279740 307770
rect 279896 305590 279924 307838
rect 279884 305584 279936 305590
rect 279884 305526 279936 305532
rect 279988 304706 280016 310420
rect 280068 309120 280120 309126
rect 280068 309062 280120 309068
rect 279976 304700 280028 304706
rect 279976 304642 280028 304648
rect 279528 302206 279740 302234
rect 279528 15910 279556 302206
rect 279976 300416 280028 300422
rect 279976 300358 280028 300364
rect 279884 244860 279936 244866
rect 279884 244802 279936 244808
rect 279896 154290 279924 244802
rect 279988 157078 280016 300358
rect 279976 157072 280028 157078
rect 279976 157014 280028 157020
rect 280080 155922 280108 309062
rect 280172 307873 280200 310420
rect 280158 307864 280214 307873
rect 280356 307834 280384 310420
rect 280158 307799 280214 307808
rect 280344 307828 280396 307834
rect 280344 307770 280396 307776
rect 280540 306354 280568 310420
rect 280724 308038 280752 310420
rect 280712 308032 280764 308038
rect 280712 307974 280764 307980
rect 280908 306354 280936 310420
rect 280988 307828 281040 307834
rect 280988 307770 281040 307776
rect 280344 306332 280396 306338
rect 280344 306274 280396 306280
rect 280448 306326 280568 306354
rect 280724 306326 280936 306354
rect 280068 155916 280120 155922
rect 280068 155858 280120 155864
rect 280080 155650 280108 155858
rect 280068 155644 280120 155650
rect 280068 155586 280120 155592
rect 279884 154284 279936 154290
rect 279884 154226 279936 154232
rect 280356 145586 280384 306274
rect 280448 152522 280476 306326
rect 280528 306196 280580 306202
rect 280528 306138 280580 306144
rect 280436 152516 280488 152522
rect 280436 152458 280488 152464
rect 280344 145580 280396 145586
rect 280344 145522 280396 145528
rect 280540 111110 280568 306138
rect 280724 134570 280752 306326
rect 281000 306218 281028 307770
rect 281092 306338 281120 310420
rect 281276 307902 281304 310420
rect 281264 307896 281316 307902
rect 281264 307838 281316 307844
rect 281080 306332 281132 306338
rect 281080 306274 281132 306280
rect 280816 306190 281028 306218
rect 281460 306202 281488 310420
rect 281448 306196 281500 306202
rect 280712 134564 280764 134570
rect 280712 134506 280764 134512
rect 280528 111104 280580 111110
rect 280528 111046 280580 111052
rect 279516 15904 279568 15910
rect 279516 15846 279568 15852
rect 280816 10334 280844 306190
rect 281448 306138 281500 306144
rect 281540 306196 281592 306202
rect 281540 306138 281592 306144
rect 280894 306096 280950 306105
rect 280894 306031 280950 306040
rect 280908 157457 280936 306031
rect 281448 305584 281500 305590
rect 281448 305526 281500 305532
rect 281264 250708 281316 250714
rect 281264 250650 281316 250656
rect 280988 193860 281040 193866
rect 280988 193802 281040 193808
rect 281000 159730 281028 193802
rect 280988 159724 281040 159730
rect 280988 159666 281040 159672
rect 281276 158982 281304 250650
rect 281356 246900 281408 246906
rect 281356 246842 281408 246848
rect 281264 158976 281316 158982
rect 281264 158918 281316 158924
rect 281368 157570 281396 246842
rect 281460 158302 281488 305526
rect 281552 305522 281580 306138
rect 281540 305516 281592 305522
rect 281540 305458 281592 305464
rect 281448 158296 281500 158302
rect 281448 158238 281500 158244
rect 281368 157542 281488 157570
rect 280894 157448 280950 157457
rect 280894 157383 280950 157392
rect 281460 155650 281488 157542
rect 281448 155644 281500 155650
rect 281448 155586 281500 155592
rect 281460 155514 281488 155586
rect 281448 155508 281500 155514
rect 281448 155450 281500 155456
rect 281644 17338 281672 310420
rect 281724 306400 281776 306406
rect 281724 306342 281776 306348
rect 281736 124914 281764 306342
rect 281828 138718 281856 310420
rect 281908 306332 281960 306338
rect 281908 306274 281960 306280
rect 281920 146946 281948 306274
rect 282012 148374 282040 310420
rect 282196 306338 282224 310420
rect 282380 306406 282408 310420
rect 282368 306400 282420 306406
rect 282368 306342 282420 306348
rect 282184 306332 282236 306338
rect 282184 306274 282236 306280
rect 282276 306332 282328 306338
rect 282276 306274 282328 306280
rect 282288 305454 282316 306274
rect 282276 305448 282328 305454
rect 282276 305390 282328 305396
rect 282564 296714 282592 310420
rect 282644 309052 282696 309058
rect 282644 308994 282696 309000
rect 282656 305674 282684 308994
rect 282748 307834 282776 310420
rect 282828 308372 282880 308378
rect 282828 308314 282880 308320
rect 282736 307828 282788 307834
rect 282736 307770 282788 307776
rect 282656 305646 282776 305674
rect 282644 303612 282696 303618
rect 282644 303554 282696 303560
rect 282104 296686 282592 296714
rect 282000 148368 282052 148374
rect 282000 148310 282052 148316
rect 282000 147008 282052 147014
rect 282000 146950 282052 146956
rect 281908 146940 281960 146946
rect 281908 146882 281960 146888
rect 281816 138712 281868 138718
rect 281816 138654 281868 138660
rect 281724 124908 281776 124914
rect 281724 124850 281776 124856
rect 281632 17332 281684 17338
rect 281632 17274 281684 17280
rect 280804 10328 280856 10334
rect 280804 10270 280856 10276
rect 282012 6914 282040 146950
rect 281920 6886 282040 6914
rect 279424 4956 279476 4962
rect 279424 4898 279476 4904
rect 280712 3188 280764 3194
rect 280712 3130 280764 3136
rect 280724 480 280752 3130
rect 281920 480 281948 6886
rect 282104 4418 282132 296686
rect 282552 248260 282604 248266
rect 282552 248202 282604 248208
rect 282564 158642 282592 248202
rect 282656 171086 282684 303554
rect 282644 171080 282696 171086
rect 282644 171022 282696 171028
rect 282656 170406 282684 171022
rect 282644 170400 282696 170406
rect 282644 170342 282696 170348
rect 282552 158636 282604 158642
rect 282552 158578 282604 158584
rect 282748 157214 282776 305646
rect 282736 157208 282788 157214
rect 282736 157150 282788 157156
rect 282748 156806 282776 157150
rect 282840 157146 282868 308314
rect 282932 306354 282960 310420
rect 283116 307873 283144 310420
rect 283102 307864 283158 307873
rect 283102 307799 283158 307808
rect 283300 306354 283328 310420
rect 282932 306326 283052 306354
rect 282920 305108 282972 305114
rect 282920 305050 282972 305056
rect 282828 157140 282880 157146
rect 282828 157082 282880 157088
rect 282736 156800 282788 156806
rect 282736 156742 282788 156748
rect 282182 125488 282238 125497
rect 282182 125423 282238 125432
rect 282092 4412 282144 4418
rect 282092 4354 282144 4360
rect 282196 3534 282224 125423
rect 282184 3528 282236 3534
rect 282184 3470 282236 3476
rect 282932 3482 282960 305050
rect 283024 3602 283052 306326
rect 283208 306326 283328 306354
rect 283104 302796 283156 302802
rect 283104 302738 283156 302744
rect 283116 6914 283144 302738
rect 283208 11626 283236 306326
rect 283484 302234 283512 310420
rect 283668 302802 283696 310420
rect 283656 302796 283708 302802
rect 283656 302738 283708 302744
rect 283300 302206 283512 302234
rect 283300 88806 283328 302206
rect 283852 296714 283880 310420
rect 284036 305114 284064 310420
rect 284116 308712 284168 308718
rect 284116 308654 284168 308660
rect 284024 305108 284076 305114
rect 284024 305050 284076 305056
rect 284128 302234 284156 308654
rect 284220 307834 284248 310420
rect 284208 307828 284260 307834
rect 284208 307770 284260 307776
rect 284404 306626 284432 310420
rect 284484 307828 284536 307834
rect 284484 307770 284536 307776
rect 284220 306598 284432 306626
rect 284220 306374 284248 306598
rect 284496 306374 284524 307770
rect 284220 306346 284340 306374
rect 284128 302206 284248 302234
rect 284116 300484 284168 300490
rect 284116 300426 284168 300432
rect 283392 296686 283880 296714
rect 283392 147014 283420 296686
rect 283932 250776 283984 250782
rect 283932 250718 283984 250724
rect 283944 248414 283972 250718
rect 283944 248386 284064 248414
rect 283932 248056 283984 248062
rect 283932 247998 283984 248004
rect 283944 247081 283972 247998
rect 283930 247072 283986 247081
rect 283930 247007 283986 247016
rect 283564 191888 283616 191894
rect 283564 191830 283616 191836
rect 283576 159798 283604 191830
rect 283564 159792 283616 159798
rect 283564 159734 283616 159740
rect 284036 158914 284064 248386
rect 284024 158908 284076 158914
rect 284024 158850 284076 158856
rect 284128 155854 284156 300426
rect 284116 155848 284168 155854
rect 284116 155790 284168 155796
rect 284220 154358 284248 302206
rect 284208 154352 284260 154358
rect 284208 154294 284260 154300
rect 283380 147008 283432 147014
rect 283380 146950 283432 146956
rect 283288 88800 283340 88806
rect 283288 88742 283340 88748
rect 283196 11620 283248 11626
rect 283196 11562 283248 11568
rect 283116 6886 283236 6914
rect 283012 3596 283064 3602
rect 283012 3538 283064 3544
rect 282932 3454 283144 3482
rect 283116 480 283144 3454
rect 283208 3194 283236 6886
rect 284312 3602 284340 306346
rect 284404 306346 284524 306374
rect 284300 3596 284352 3602
rect 284300 3538 284352 3544
rect 284404 3482 284432 306346
rect 284588 306218 284616 310420
rect 284668 306400 284720 306406
rect 284668 306342 284720 306348
rect 284312 3454 284432 3482
rect 284496 306190 284616 306218
rect 283196 3188 283248 3194
rect 283196 3130 283248 3136
rect 284312 480 284340 3454
rect 284496 3058 284524 306190
rect 284576 305516 284628 305522
rect 284576 305458 284628 305464
rect 284588 6934 284616 305458
rect 284680 8974 284708 306342
rect 284772 154630 284800 310420
rect 284956 305522 284984 310420
rect 285036 308848 285088 308854
rect 285036 308790 285088 308796
rect 284944 305516 284996 305522
rect 284944 305458 284996 305464
rect 285048 296714 285076 308790
rect 285140 307902 285168 310420
rect 285128 307896 285180 307902
rect 285128 307838 285180 307844
rect 285324 307834 285352 310420
rect 285312 307828 285364 307834
rect 285312 307770 285364 307776
rect 285508 306406 285536 310420
rect 285692 306542 285720 310420
rect 285876 309134 285904 310420
rect 285784 309106 285904 309134
rect 285680 306536 285732 306542
rect 285680 306478 285732 306484
rect 285496 306400 285548 306406
rect 285496 306342 285548 306348
rect 285680 306400 285732 306406
rect 285680 306342 285732 306348
rect 285496 302796 285548 302802
rect 285496 302738 285548 302744
rect 285404 300552 285456 300558
rect 285404 300494 285456 300500
rect 284956 296686 285076 296714
rect 284956 158846 284984 296686
rect 285036 247784 285088 247790
rect 285036 247726 285088 247732
rect 285048 247081 285076 247726
rect 285034 247072 285090 247081
rect 285034 247007 285090 247016
rect 284944 158840 284996 158846
rect 284944 158782 284996 158788
rect 285416 158234 285444 300494
rect 285404 158228 285456 158234
rect 285404 158170 285456 158176
rect 285508 158098 285536 302738
rect 285588 246356 285640 246362
rect 285588 246298 285640 246304
rect 285496 158092 285548 158098
rect 285496 158034 285548 158040
rect 284760 154624 284812 154630
rect 284760 154566 284812 154572
rect 284668 8968 284720 8974
rect 284668 8910 284720 8916
rect 284576 6928 284628 6934
rect 284576 6870 284628 6876
rect 285600 4146 285628 246298
rect 285692 5098 285720 306342
rect 285784 6526 285812 309106
rect 286060 308106 286088 310420
rect 286048 308100 286100 308106
rect 286048 308042 286100 308048
rect 286244 307970 286272 310420
rect 286232 307964 286284 307970
rect 286232 307906 286284 307912
rect 286324 307828 286376 307834
rect 286324 307770 286376 307776
rect 286048 306536 286100 306542
rect 286048 306478 286100 306484
rect 286140 306536 286192 306542
rect 286140 306478 286192 306484
rect 285956 306400 286008 306406
rect 285956 306342 286008 306348
rect 285864 305516 285916 305522
rect 285864 305458 285916 305464
rect 285876 148374 285904 305458
rect 285968 151162 285996 306342
rect 286060 153950 286088 306478
rect 286152 159662 286180 306478
rect 286140 159656 286192 159662
rect 286140 159598 286192 159604
rect 286140 158568 286192 158574
rect 286140 158510 286192 158516
rect 286152 157962 286180 158510
rect 286140 157956 286192 157962
rect 286140 157898 286192 157904
rect 286048 153944 286100 153950
rect 286048 153886 286100 153892
rect 285956 151156 286008 151162
rect 285956 151098 286008 151104
rect 285864 148368 285916 148374
rect 285864 148310 285916 148316
rect 286336 142934 286364 307770
rect 286428 306474 286456 310420
rect 286612 306542 286640 310420
rect 286600 306536 286652 306542
rect 286600 306478 286652 306484
rect 286416 306468 286468 306474
rect 286416 306410 286468 306416
rect 286796 306406 286824 310420
rect 286784 306400 286836 306406
rect 286784 306342 286836 306348
rect 286980 305522 287008 310420
rect 287060 306400 287112 306406
rect 287060 306342 287112 306348
rect 286968 305516 287020 305522
rect 286968 305458 287020 305464
rect 286692 302864 286744 302870
rect 286692 302806 286744 302812
rect 286600 247988 286652 247994
rect 286600 247930 286652 247936
rect 286612 247081 286640 247930
rect 286598 247072 286654 247081
rect 286598 247007 286654 247016
rect 286704 158574 286732 302806
rect 286876 300620 286928 300626
rect 286876 300562 286928 300568
rect 286784 243568 286836 243574
rect 286784 243510 286836 243516
rect 286796 158574 286824 243510
rect 286692 158568 286744 158574
rect 286692 158510 286744 158516
rect 286784 158568 286836 158574
rect 286784 158510 286836 158516
rect 286888 157214 286916 300562
rect 286966 158808 287022 158817
rect 286966 158743 287022 158752
rect 286876 157208 286928 157214
rect 286876 157150 286928 157156
rect 286324 142928 286376 142934
rect 286324 142870 286376 142876
rect 285772 6520 285824 6526
rect 285772 6462 285824 6468
rect 286980 6390 287008 158743
rect 287072 51746 287100 306342
rect 287164 305522 287192 310420
rect 287348 306354 287376 310420
rect 287256 306326 287376 306354
rect 287152 305516 287204 305522
rect 287152 305458 287204 305464
rect 287152 305380 287204 305386
rect 287152 305322 287204 305328
rect 287164 134570 287192 305322
rect 287256 146946 287284 306326
rect 287532 306218 287560 310420
rect 287612 309120 287664 309126
rect 287612 309062 287664 309068
rect 287624 308786 287652 309062
rect 287612 308780 287664 308786
rect 287612 308722 287664 308728
rect 287348 306190 287560 306218
rect 287348 153882 287376 306190
rect 287716 306082 287744 310420
rect 287796 307896 287848 307902
rect 287796 307838 287848 307844
rect 287440 306054 287744 306082
rect 287440 156738 287468 306054
rect 287520 305516 287572 305522
rect 287520 305458 287572 305464
rect 287532 159594 287560 305458
rect 287808 296714 287836 307838
rect 287900 306406 287928 310420
rect 287888 306400 287940 306406
rect 287888 306342 287940 306348
rect 288084 305386 288112 310420
rect 288268 307873 288296 310420
rect 288254 307864 288310 307873
rect 288254 307799 288310 307808
rect 288452 305522 288480 310420
rect 288636 306354 288664 310420
rect 288820 307834 288848 310420
rect 288808 307828 288860 307834
rect 288808 307770 288860 307776
rect 288544 306326 288664 306354
rect 288716 306400 288768 306406
rect 289004 306354 289032 310420
rect 288716 306342 288768 306348
rect 288440 305516 288492 305522
rect 288440 305458 288492 305464
rect 288072 305380 288124 305386
rect 288072 305322 288124 305328
rect 288440 305380 288492 305386
rect 288440 305322 288492 305328
rect 288072 300688 288124 300694
rect 288072 300630 288124 300636
rect 287716 296686 287836 296714
rect 287520 159588 287572 159594
rect 287520 159530 287572 159536
rect 287428 156732 287480 156738
rect 287428 156674 287480 156680
rect 287428 154624 287480 154630
rect 287428 154566 287480 154572
rect 287336 153876 287388 153882
rect 287336 153818 287388 153824
rect 287244 146940 287296 146946
rect 287244 146882 287296 146888
rect 287152 134564 287204 134570
rect 287152 134506 287204 134512
rect 287060 51740 287112 51746
rect 287060 51682 287112 51688
rect 286968 6384 287020 6390
rect 286968 6326 287020 6332
rect 285680 5092 285732 5098
rect 285680 5034 285732 5040
rect 285588 4140 285640 4146
rect 285588 4082 285640 4088
rect 285036 3596 285088 3602
rect 285036 3538 285088 3544
rect 284484 3052 284536 3058
rect 284484 2994 284536 3000
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285048 354 285076 3538
rect 286600 3052 286652 3058
rect 286600 2994 286652 3000
rect 286612 480 286640 2994
rect 285374 354 285486 480
rect 285048 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287440 354 287468 154566
rect 287716 4214 287744 296686
rect 287796 247920 287848 247926
rect 287796 247862 287848 247868
rect 287808 247081 287836 247862
rect 287794 247072 287850 247081
rect 287794 247007 287850 247016
rect 288084 158710 288112 300630
rect 288348 251184 288400 251190
rect 288348 251126 288400 251132
rect 288256 247444 288308 247450
rect 288256 247386 288308 247392
rect 288164 244656 288216 244662
rect 288164 244598 288216 244604
rect 288176 244361 288204 244598
rect 288162 244352 288218 244361
rect 288162 244287 288218 244296
rect 288268 243114 288296 247386
rect 288176 243086 288296 243114
rect 288072 158704 288124 158710
rect 288072 158646 288124 158652
rect 288176 158506 288204 243086
rect 288360 238754 288388 251126
rect 288268 238726 288388 238754
rect 288268 159526 288296 238726
rect 288256 159520 288308 159526
rect 288256 159462 288308 159468
rect 288346 158808 288402 158817
rect 288346 158743 288402 158752
rect 288256 158704 288308 158710
rect 288256 158646 288308 158652
rect 288164 158500 288216 158506
rect 288164 158442 288216 158448
rect 288268 157894 288296 158646
rect 288256 157888 288308 157894
rect 288256 157830 288308 157836
rect 288360 6186 288388 158743
rect 288452 6866 288480 305322
rect 288544 14482 288572 306326
rect 288624 305448 288676 305454
rect 288624 305390 288676 305396
rect 288636 133210 288664 305390
rect 288728 145586 288756 306342
rect 288820 306326 289032 306354
rect 288820 149802 288848 306326
rect 288900 305516 288952 305522
rect 288900 305458 288952 305464
rect 288912 152726 288940 305458
rect 289188 305386 289216 310420
rect 289176 305380 289228 305386
rect 289176 305322 289228 305328
rect 289372 302234 289400 310420
rect 289450 308952 289506 308961
rect 289450 308887 289506 308896
rect 289004 302206 289400 302234
rect 289004 159905 289032 302206
rect 289464 296714 289492 308887
rect 289556 306406 289584 310420
rect 289544 306400 289596 306406
rect 289544 306342 289596 306348
rect 289740 305454 289768 310420
rect 289820 306536 289872 306542
rect 289820 306478 289872 306484
rect 289728 305448 289780 305454
rect 289728 305390 289780 305396
rect 289544 300756 289596 300762
rect 289544 300698 289596 300704
rect 289096 296686 289492 296714
rect 288990 159896 289046 159905
rect 288990 159831 289046 159840
rect 289096 158778 289124 296686
rect 289176 247852 289228 247858
rect 289176 247794 289228 247800
rect 289188 247081 289216 247794
rect 289174 247072 289230 247081
rect 289174 247007 289230 247016
rect 289084 158772 289136 158778
rect 289084 158714 289136 158720
rect 289556 158030 289584 300698
rect 289636 250368 289688 250374
rect 289636 250310 289688 250316
rect 289648 159458 289676 250310
rect 289636 159452 289688 159458
rect 289636 159394 289688 159400
rect 289726 158808 289782 158817
rect 289726 158743 289782 158752
rect 289360 158024 289412 158030
rect 289360 157966 289412 157972
rect 289544 158024 289596 158030
rect 289544 157966 289596 157972
rect 289372 157622 289400 157966
rect 289360 157616 289412 157622
rect 289360 157558 289412 157564
rect 288900 152720 288952 152726
rect 288900 152662 288952 152668
rect 288808 149796 288860 149802
rect 288808 149738 288860 149744
rect 288716 145580 288768 145586
rect 288716 145522 288768 145528
rect 288624 133204 288676 133210
rect 288624 133146 288676 133152
rect 288532 14476 288584 14482
rect 288532 14418 288584 14424
rect 288992 6928 289044 6934
rect 288992 6870 289044 6876
rect 288440 6860 288492 6866
rect 288440 6802 288492 6808
rect 288348 6180 288400 6186
rect 288348 6122 288400 6128
rect 287704 4208 287756 4214
rect 287704 4150 287756 4156
rect 289004 480 289032 6870
rect 289740 6254 289768 158743
rect 289728 6248 289780 6254
rect 289728 6190 289780 6196
rect 289832 5166 289860 306478
rect 289924 306474 289952 310420
rect 289912 306468 289964 306474
rect 289912 306410 289964 306416
rect 290108 306354 290136 310420
rect 290016 306326 290136 306354
rect 290188 306400 290240 306406
rect 290188 306342 290240 306348
rect 289912 305448 289964 305454
rect 289912 305390 289964 305396
rect 289820 5160 289872 5166
rect 289820 5102 289872 5108
rect 289924 5030 289952 305390
rect 290016 6798 290044 306326
rect 290096 305516 290148 305522
rect 290096 305458 290148 305464
rect 290108 22778 290136 305458
rect 290200 89010 290228 306342
rect 290292 89078 290320 310420
rect 290372 306468 290424 306474
rect 290372 306410 290424 306416
rect 290384 244769 290412 306410
rect 290476 305454 290504 310420
rect 290660 305522 290688 310420
rect 290740 308032 290792 308038
rect 290740 307974 290792 307980
rect 290648 305516 290700 305522
rect 290648 305458 290700 305464
rect 290464 305448 290516 305454
rect 290464 305390 290516 305396
rect 290370 244760 290426 244769
rect 290370 244695 290426 244704
rect 290646 158808 290702 158817
rect 290646 158743 290702 158752
rect 290280 89072 290332 89078
rect 290280 89014 290332 89020
rect 290188 89004 290240 89010
rect 290188 88946 290240 88952
rect 290096 22772 290148 22778
rect 290096 22714 290148 22720
rect 290004 6792 290056 6798
rect 290004 6734 290056 6740
rect 290660 6458 290688 158743
rect 290752 157350 290780 307974
rect 290844 306406 290872 310420
rect 291028 306542 291056 310420
rect 291016 306536 291068 306542
rect 291016 306478 291068 306484
rect 291212 306474 291240 310420
rect 291396 309134 291424 310420
rect 291304 309106 291424 309134
rect 291200 306468 291252 306474
rect 291200 306410 291252 306416
rect 290832 306400 290884 306406
rect 290832 306342 290884 306348
rect 291304 305504 291332 309106
rect 291476 306468 291528 306474
rect 291476 306410 291528 306416
rect 291212 305476 291332 305504
rect 291384 305516 291436 305522
rect 290924 250980 290976 250986
rect 290924 250922 290976 250928
rect 290832 245472 290884 245478
rect 290832 245414 290884 245420
rect 290844 244497 290872 245414
rect 290830 244488 290886 244497
rect 290830 244423 290886 244432
rect 290832 243704 290884 243710
rect 290832 243646 290884 243652
rect 290844 158710 290872 243646
rect 290936 159254 290964 250922
rect 291016 250912 291068 250918
rect 291016 250854 291068 250860
rect 291028 159322 291056 250854
rect 291108 245064 291160 245070
rect 291108 245006 291160 245012
rect 291120 244361 291148 245006
rect 291106 244352 291162 244361
rect 291106 244287 291162 244296
rect 291016 159316 291068 159322
rect 291016 159258 291068 159264
rect 290924 159248 290976 159254
rect 290924 159190 290976 159196
rect 291106 158808 291162 158817
rect 291106 158743 291162 158752
rect 290832 158704 290884 158710
rect 290832 158646 290884 158652
rect 290740 157344 290792 157350
rect 290740 157286 290792 157292
rect 290752 156602 290780 157286
rect 290740 156596 290792 156602
rect 290740 156538 290792 156544
rect 290648 6452 290700 6458
rect 290648 6394 290700 6400
rect 289912 5024 289964 5030
rect 289912 4966 289964 4972
rect 290188 4208 290240 4214
rect 290188 4150 290240 4156
rect 290200 480 290228 4150
rect 291120 3670 291148 158743
rect 291212 18630 291240 305476
rect 291384 305458 291436 305464
rect 291292 305380 291344 305386
rect 291292 305322 291344 305328
rect 291304 141438 291332 305322
rect 291396 142866 291424 305458
rect 291488 144226 291516 306410
rect 291580 306354 291608 310420
rect 291580 306326 291700 306354
rect 291568 305448 291620 305454
rect 291568 305390 291620 305396
rect 291580 151094 291608 305390
rect 291672 152658 291700 306326
rect 291764 305522 291792 310420
rect 291948 308106 291976 310420
rect 291844 308100 291896 308106
rect 291844 308042 291896 308048
rect 291936 308100 291988 308106
rect 291936 308042 291988 308048
rect 291752 305516 291804 305522
rect 291752 305458 291804 305464
rect 291752 244384 291804 244390
rect 291750 244352 291752 244361
rect 291804 244352 291806 244361
rect 291750 244287 291806 244296
rect 291660 152652 291712 152658
rect 291660 152594 291712 152600
rect 291568 151088 291620 151094
rect 291568 151030 291620 151036
rect 291476 144220 291528 144226
rect 291476 144162 291528 144168
rect 291476 142928 291528 142934
rect 291476 142870 291528 142876
rect 291384 142860 291436 142866
rect 291384 142802 291436 142808
rect 291292 141432 291344 141438
rect 291292 141374 291344 141380
rect 291200 18624 291252 18630
rect 291200 18566 291252 18572
rect 291488 6914 291516 142870
rect 291396 6886 291516 6914
rect 291108 3664 291160 3670
rect 291108 3606 291160 3612
rect 291396 480 291424 6886
rect 291856 3534 291884 308042
rect 291936 307828 291988 307834
rect 291936 307770 291988 307776
rect 291948 156670 291976 307770
rect 292132 305454 292160 310420
rect 292120 305448 292172 305454
rect 292120 305390 292172 305396
rect 292316 305386 292344 310420
rect 292500 308689 292528 310420
rect 292486 308680 292542 308689
rect 292486 308615 292542 308624
rect 292684 306592 292712 310420
rect 292500 306564 292712 306592
rect 292396 305516 292448 305522
rect 292396 305458 292448 305464
rect 292304 305380 292356 305386
rect 292304 305322 292356 305328
rect 292408 302234 292436 305458
rect 292500 304298 292528 306564
rect 292672 306468 292724 306474
rect 292672 306410 292724 306416
rect 292580 306400 292632 306406
rect 292580 306342 292632 306348
rect 292488 304292 292540 304298
rect 292488 304234 292540 304240
rect 292316 302206 292436 302234
rect 292120 245404 292172 245410
rect 292120 245346 292172 245352
rect 292132 244361 292160 245346
rect 292118 244352 292174 244361
rect 292118 244287 292174 244296
rect 292316 158438 292344 302206
rect 292396 251048 292448 251054
rect 292396 250990 292448 250996
rect 292408 158846 292436 250990
rect 292396 158840 292448 158846
rect 292396 158782 292448 158788
rect 292486 158808 292542 158817
rect 292486 158743 292542 158752
rect 292304 158432 292356 158438
rect 292304 158374 292356 158380
rect 292316 158166 292344 158374
rect 292304 158160 292356 158166
rect 292304 158102 292356 158108
rect 292394 157448 292450 157457
rect 292394 157383 292450 157392
rect 291936 156664 291988 156670
rect 291936 156606 291988 156612
rect 292408 16574 292436 157383
rect 292316 16546 292436 16574
rect 291844 3528 291896 3534
rect 291844 3470 291896 3476
rect 292316 3466 292344 16546
rect 292500 11778 292528 158743
rect 292592 130422 292620 306342
rect 292684 138718 292712 306410
rect 292868 306354 292896 310420
rect 292948 306536 293000 306542
rect 292948 306478 293000 306484
rect 292776 306326 292896 306354
rect 292776 140078 292804 306326
rect 292960 304450 292988 306478
rect 293052 306406 293080 310420
rect 293236 306542 293264 310420
rect 293316 307964 293368 307970
rect 293316 307906 293368 307912
rect 293224 306536 293276 306542
rect 293224 306478 293276 306484
rect 293040 306400 293092 306406
rect 293040 306342 293092 306348
rect 293328 306082 293356 307906
rect 293420 306474 293448 310420
rect 293500 308100 293552 308106
rect 293500 308042 293552 308048
rect 293408 306468 293460 306474
rect 293408 306410 293460 306416
rect 292868 304422 292988 304450
rect 293236 306054 293356 306082
rect 292868 149734 292896 304422
rect 292948 304292 293000 304298
rect 292948 304234 293000 304240
rect 292960 246362 292988 304234
rect 292948 246356 293000 246362
rect 292948 246298 293000 246304
rect 292948 153944 293000 153950
rect 292948 153886 293000 153892
rect 292856 149728 292908 149734
rect 292856 149670 292908 149676
rect 292764 140072 292816 140078
rect 292764 140014 292816 140020
rect 292672 138712 292724 138718
rect 292672 138654 292724 138660
rect 292580 130416 292632 130422
rect 292580 130358 292632 130364
rect 292960 12434 292988 153886
rect 293236 16574 293264 306054
rect 293512 302234 293540 308042
rect 293604 307834 293632 310420
rect 293788 307873 293816 310420
rect 293774 307864 293830 307873
rect 293592 307828 293644 307834
rect 293774 307799 293830 307808
rect 293592 307770 293644 307776
rect 293972 306474 294000 310420
rect 293960 306468 294012 306474
rect 293960 306410 294012 306416
rect 294052 306400 294104 306406
rect 293972 306348 294052 306354
rect 293972 306342 294104 306348
rect 293972 306326 294092 306342
rect 293684 302728 293736 302734
rect 293684 302670 293736 302676
rect 293328 302206 293540 302234
rect 293328 131782 293356 302206
rect 293592 251116 293644 251122
rect 293592 251058 293644 251064
rect 293408 248396 293460 248402
rect 293408 248338 293460 248344
rect 293420 247081 293448 248338
rect 293500 247580 293552 247586
rect 293500 247522 293552 247528
rect 293406 247072 293462 247081
rect 293406 247007 293462 247016
rect 293408 244928 293460 244934
rect 293408 244870 293460 244876
rect 293420 244769 293448 244870
rect 293406 244760 293462 244769
rect 293406 244695 293462 244704
rect 293512 239834 293540 247522
rect 293500 239828 293552 239834
rect 293500 239770 293552 239776
rect 293604 159186 293632 251058
rect 293592 159180 293644 159186
rect 293592 159122 293644 159128
rect 293498 158808 293554 158817
rect 293498 158743 293554 158752
rect 293316 131776 293368 131782
rect 293316 131718 293368 131724
rect 293236 16546 293356 16574
rect 292960 12406 293264 12434
rect 292408 11750 292528 11778
rect 292408 4078 292436 11750
rect 292488 8968 292540 8974
rect 292488 8910 292540 8916
rect 292396 4072 292448 4078
rect 292396 4014 292448 4020
rect 292500 3482 292528 8910
rect 292304 3460 292356 3466
rect 292500 3454 292620 3482
rect 292304 3402 292356 3408
rect 292592 480 292620 3454
rect 287766 354 287878 480
rect 287440 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 12406
rect 293328 5506 293356 16546
rect 293316 5500 293368 5506
rect 293316 5442 293368 5448
rect 293512 3330 293540 158743
rect 293696 158438 293724 302670
rect 293776 245336 293828 245342
rect 293774 245304 293776 245313
rect 293828 245304 293830 245313
rect 293774 245239 293830 245248
rect 293774 245168 293830 245177
rect 293774 245103 293830 245112
rect 293788 244361 293816 245103
rect 293868 244520 293920 244526
rect 293868 244462 293920 244468
rect 293774 244352 293830 244361
rect 293774 244287 293830 244296
rect 293776 239828 293828 239834
rect 293776 239770 293828 239776
rect 293788 168366 293816 239770
rect 293776 168360 293828 168366
rect 293776 168302 293828 168308
rect 293774 167104 293830 167113
rect 293774 167039 293830 167048
rect 293684 158432 293736 158438
rect 293684 158374 293736 158380
rect 293590 149152 293646 149161
rect 293590 149087 293646 149096
rect 293604 6322 293632 149087
rect 293592 6316 293644 6322
rect 293592 6258 293644 6264
rect 293788 3874 293816 167039
rect 293880 3942 293908 244462
rect 293972 4894 294000 306326
rect 294052 305448 294104 305454
rect 294052 305390 294104 305396
rect 294064 6662 294092 305390
rect 294156 305232 294184 310420
rect 294340 306406 294368 310420
rect 294328 306400 294380 306406
rect 294328 306342 294380 306348
rect 294156 305204 294276 305232
rect 294144 305108 294196 305114
rect 294144 305050 294196 305056
rect 294156 6730 294184 305050
rect 294248 9178 294276 305204
rect 294524 305114 294552 310420
rect 294708 307902 294736 310420
rect 294696 307896 294748 307902
rect 294696 307838 294748 307844
rect 294604 307828 294656 307834
rect 294604 307770 294656 307776
rect 294512 305108 294564 305114
rect 294512 305050 294564 305056
rect 294616 304994 294644 307770
rect 294432 304966 294644 304994
rect 294432 302258 294460 304966
rect 294892 304858 294920 310420
rect 294972 309120 295024 309126
rect 294972 309062 295024 309068
rect 294524 304830 294920 304858
rect 294420 302252 294472 302258
rect 294420 302194 294472 302200
rect 294524 296714 294552 304830
rect 294604 302252 294656 302258
rect 294604 302194 294656 302200
rect 294340 296686 294552 296714
rect 294340 159769 294368 296686
rect 294326 159760 294382 159769
rect 294326 159695 294382 159704
rect 294328 155712 294380 155718
rect 294328 155654 294380 155660
rect 294340 154902 294368 155654
rect 294328 154896 294380 154902
rect 294328 154838 294380 154844
rect 294616 9246 294644 302194
rect 294984 296714 295012 309062
rect 295076 305454 295104 310420
rect 295260 307834 295288 310420
rect 295444 307970 295472 310420
rect 295432 307964 295484 307970
rect 295432 307906 295484 307912
rect 295248 307828 295300 307834
rect 295248 307770 295300 307776
rect 295340 306400 295392 306406
rect 295628 306354 295656 310420
rect 295340 306342 295392 306348
rect 295064 305448 295116 305454
rect 295064 305390 295116 305396
rect 294708 296686 295012 296714
rect 294708 159390 294736 296686
rect 295064 247104 295116 247110
rect 295062 247072 295064 247081
rect 295116 247072 295118 247081
rect 295062 247007 295118 247016
rect 295156 247036 295208 247042
rect 295156 246978 295208 246984
rect 294972 243636 295024 243642
rect 294972 243578 295024 243584
rect 294878 195256 294934 195265
rect 294878 195191 294934 195200
rect 294696 159384 294748 159390
rect 294696 159326 294748 159332
rect 294892 16574 294920 195191
rect 294984 155718 295012 243578
rect 295168 195974 295196 246978
rect 295248 245540 295300 245546
rect 295248 245482 295300 245488
rect 295260 244905 295288 245482
rect 295246 244896 295302 244905
rect 295246 244831 295302 244840
rect 295248 244656 295300 244662
rect 295248 244598 295300 244604
rect 295156 195968 295208 195974
rect 295156 195910 295208 195916
rect 295062 158808 295118 158817
rect 295062 158743 295118 158752
rect 294972 155712 295024 155718
rect 294972 155654 295024 155660
rect 294892 16546 295012 16574
rect 294604 9240 294656 9246
rect 294604 9182 294656 9188
rect 294236 9172 294288 9178
rect 294236 9114 294288 9120
rect 294144 6724 294196 6730
rect 294144 6666 294196 6672
rect 294052 6656 294104 6662
rect 294052 6598 294104 6604
rect 294880 6520 294932 6526
rect 294880 6462 294932 6468
rect 293960 4888 294012 4894
rect 293960 4830 294012 4836
rect 293868 3936 293920 3942
rect 293868 3878 293920 3884
rect 293776 3868 293828 3874
rect 293776 3810 293828 3816
rect 293500 3324 293552 3330
rect 293500 3266 293552 3272
rect 294892 480 294920 6462
rect 294984 3806 295012 16546
rect 295076 8974 295104 158743
rect 295064 8968 295116 8974
rect 295064 8910 295116 8916
rect 295260 4010 295288 244598
rect 295352 4826 295380 306342
rect 295444 306326 295656 306354
rect 295444 6594 295472 306326
rect 295524 305448 295576 305454
rect 295524 305390 295576 305396
rect 295536 7682 295564 305390
rect 295812 296714 295840 310420
rect 295892 306468 295944 306474
rect 295892 306410 295944 306416
rect 295904 302234 295932 306410
rect 295996 306406 296024 310420
rect 296076 307828 296128 307834
rect 296076 307770 296128 307776
rect 295984 306400 296036 306406
rect 295984 306342 296036 306348
rect 295904 302206 296024 302234
rect 295628 296686 295840 296714
rect 295628 152590 295656 296686
rect 295798 245440 295854 245449
rect 295798 245375 295854 245384
rect 295812 244905 295840 245375
rect 295798 244896 295854 244905
rect 295798 244831 295854 244840
rect 295708 157344 295760 157350
rect 295708 157286 295760 157292
rect 295720 156398 295748 157286
rect 295708 156392 295760 156398
rect 295708 156334 295760 156340
rect 295708 155508 295760 155514
rect 295708 155450 295760 155456
rect 295720 154970 295748 155450
rect 295708 154964 295760 154970
rect 295708 154906 295760 154912
rect 295616 152584 295668 152590
rect 295616 152526 295668 152532
rect 295524 7676 295576 7682
rect 295524 7618 295576 7624
rect 295432 6588 295484 6594
rect 295432 6530 295484 6536
rect 295340 4820 295392 4826
rect 295340 4762 295392 4768
rect 295248 4004 295300 4010
rect 295248 3946 295300 3952
rect 294972 3800 295024 3806
rect 294972 3742 295024 3748
rect 295996 3398 296024 302206
rect 296088 9110 296116 307770
rect 296180 305454 296208 310420
rect 296260 307896 296312 307902
rect 296364 307873 296392 310420
rect 296548 307873 296576 310420
rect 296260 307838 296312 307844
rect 296350 307864 296406 307873
rect 296168 305448 296220 305454
rect 296168 305390 296220 305396
rect 296272 302234 296300 307838
rect 296350 307799 296406 307808
rect 296534 307864 296590 307873
rect 296534 307799 296590 307808
rect 296732 306610 296760 310420
rect 296720 306604 296772 306610
rect 296720 306546 296772 306552
rect 296916 306490 296944 310420
rect 296732 306462 296944 306490
rect 296536 305176 296588 305182
rect 296536 305118 296588 305124
rect 296180 302206 296300 302234
rect 296180 129062 296208 302206
rect 296444 250436 296496 250442
rect 296444 250378 296496 250384
rect 296352 247648 296404 247654
rect 296352 247590 296404 247596
rect 296364 157350 296392 247590
rect 296456 159050 296484 250378
rect 296444 159044 296496 159050
rect 296444 158986 296496 158992
rect 296352 157344 296404 157350
rect 296352 157286 296404 157292
rect 296548 155514 296576 305118
rect 296628 245200 296680 245206
rect 296628 245142 296680 245148
rect 296640 244769 296668 245142
rect 296626 244760 296682 244769
rect 296626 244695 296682 244704
rect 296626 158808 296682 158817
rect 296626 158743 296682 158752
rect 296536 155508 296588 155514
rect 296536 155450 296588 155456
rect 296168 129056 296220 129062
rect 296168 128998 296220 129004
rect 296076 9104 296128 9110
rect 296076 9046 296128 9052
rect 296640 3738 296668 158743
rect 296732 6526 296760 306462
rect 297100 306354 297128 310420
rect 297284 308689 297312 310420
rect 297270 308680 297326 308689
rect 297270 308615 297326 308624
rect 297272 307964 297324 307970
rect 297272 307906 297324 307912
rect 297180 306604 297232 306610
rect 297180 306546 297232 306552
rect 296916 306326 297128 306354
rect 296812 304972 296864 304978
rect 296812 304914 296864 304920
rect 296824 245614 296852 304914
rect 296916 249490 296944 306326
rect 297192 306218 297220 306546
rect 297100 306190 297220 306218
rect 296996 305448 297048 305454
rect 296996 305390 297048 305396
rect 296904 249484 296956 249490
rect 296904 249426 296956 249432
rect 297008 249370 297036 305390
rect 296916 249342 297036 249370
rect 296916 247761 296944 249342
rect 297100 249234 297128 306190
rect 297284 302234 297312 307906
rect 297468 304978 297496 310420
rect 297652 305454 297680 310420
rect 297836 307873 297864 310420
rect 298020 308145 298048 310420
rect 298006 308136 298062 308145
rect 298006 308071 298062 308080
rect 297822 307864 297878 307873
rect 297822 307799 297878 307808
rect 298204 306474 298232 310420
rect 298388 309134 298416 310420
rect 298296 309106 298416 309134
rect 298192 306468 298244 306474
rect 298192 306410 298244 306416
rect 298100 306400 298152 306406
rect 298100 306342 298152 306348
rect 297640 305448 297692 305454
rect 297640 305390 297692 305396
rect 297456 304972 297508 304978
rect 297456 304914 297508 304920
rect 297008 249206 297128 249234
rect 297192 302206 297312 302234
rect 297008 248033 297036 249206
rect 297192 249150 297220 302206
rect 297916 256148 297968 256154
rect 297916 256090 297968 256096
rect 297640 256080 297692 256086
rect 297640 256022 297692 256028
rect 297272 256012 297324 256018
rect 297272 255954 297324 255960
rect 297180 249144 297232 249150
rect 297180 249086 297232 249092
rect 297284 248962 297312 255954
rect 297364 249484 297416 249490
rect 297364 249426 297416 249432
rect 297100 248934 297312 248962
rect 296994 248024 297050 248033
rect 296994 247959 297050 247968
rect 296902 247752 296958 247761
rect 296902 247687 296958 247696
rect 296812 245608 296864 245614
rect 296812 245550 296864 245556
rect 297100 243506 297128 248934
rect 297180 248872 297232 248878
rect 297180 248814 297232 248820
rect 297192 245177 297220 248814
rect 297272 247512 297324 247518
rect 297272 247454 297324 247460
rect 297178 245168 297234 245177
rect 297178 245103 297234 245112
rect 297088 243500 297140 243506
rect 297088 243442 297140 243448
rect 297100 238754 297128 243442
rect 297284 243166 297312 247454
rect 297376 245041 297404 249426
rect 297456 246220 297508 246226
rect 297456 246162 297508 246168
rect 297362 245032 297418 245041
rect 297362 244967 297418 244976
rect 297362 244488 297418 244497
rect 297362 244423 297418 244432
rect 297376 244390 297404 244423
rect 297364 244384 297416 244390
rect 297364 244326 297416 244332
rect 297364 243432 297416 243438
rect 297364 243374 297416 243380
rect 297272 243160 297324 243166
rect 297272 243102 297324 243108
rect 297100 238726 297312 238754
rect 297284 196897 297312 238726
rect 297270 196888 297326 196897
rect 297270 196823 297326 196832
rect 297180 196036 297232 196042
rect 297180 195978 297232 195984
rect 297192 170610 297220 195978
rect 297272 195968 297324 195974
rect 297376 195945 297404 243374
rect 297272 195910 297324 195916
rect 297362 195936 297418 195945
rect 297284 189922 297312 195910
rect 297362 195871 297418 195880
rect 297468 193866 297496 246162
rect 297548 244792 297600 244798
rect 297548 244734 297600 244740
rect 297560 243438 297588 244734
rect 297548 243432 297600 243438
rect 297548 243374 297600 243380
rect 297548 243160 297600 243166
rect 297548 243102 297600 243108
rect 297456 193860 297508 193866
rect 297456 193802 297508 193808
rect 297468 193769 297496 193802
rect 297454 193760 297510 193769
rect 297454 193695 297510 193704
rect 297560 191049 297588 243102
rect 297546 191040 297602 191049
rect 297546 190975 297602 190984
rect 297560 190454 297588 190975
rect 297468 190426 297588 190454
rect 297272 189916 297324 189922
rect 297272 189858 297324 189864
rect 297362 189136 297418 189145
rect 297362 189071 297418 189080
rect 297180 170604 297232 170610
rect 297180 170546 297232 170552
rect 297376 157690 297404 189071
rect 297468 159866 297496 190426
rect 297652 189961 297680 256022
rect 297732 244588 297784 244594
rect 297732 244530 297784 244536
rect 297638 189952 297694 189961
rect 297638 189887 297694 189896
rect 297652 189145 297680 189887
rect 297638 189136 297694 189145
rect 297638 189071 297694 189080
rect 297546 188184 297602 188193
rect 297546 188119 297602 188128
rect 297560 159934 297588 188119
rect 297640 171080 297692 171086
rect 297640 171022 297692 171028
rect 297652 169969 297680 171022
rect 297638 169960 297694 169969
rect 297638 169895 297694 169904
rect 297640 168360 297692 168366
rect 297640 168302 297692 168308
rect 297548 159928 297600 159934
rect 297548 159870 297600 159876
rect 297456 159860 297508 159866
rect 297456 159802 297508 159808
rect 297652 159390 297680 168302
rect 297744 168065 297772 244530
rect 297824 243840 297876 243846
rect 297824 243782 297876 243788
rect 297730 168056 297786 168065
rect 297730 167991 297786 168000
rect 297640 159384 297692 159390
rect 297640 159326 297692 159332
rect 297836 158778 297864 243782
rect 297928 168337 297956 256090
rect 298008 246288 298060 246294
rect 298008 246230 298060 246236
rect 297914 168328 297970 168337
rect 297914 168263 297970 168272
rect 297928 167686 297956 168263
rect 297916 167680 297968 167686
rect 297916 167622 297968 167628
rect 297824 158772 297876 158778
rect 297824 158714 297876 158720
rect 297364 157684 297416 157690
rect 297364 157626 297416 157632
rect 298020 154494 298048 246230
rect 298008 154488 298060 154494
rect 298008 154430 298060 154436
rect 298112 10334 298140 306342
rect 298296 305368 298324 309106
rect 298468 306468 298520 306474
rect 298468 306410 298520 306416
rect 298376 305448 298428 305454
rect 298376 305390 298428 305396
rect 298204 305340 298324 305368
rect 298204 152522 298232 305340
rect 298284 305244 298336 305250
rect 298284 305186 298336 305192
rect 298296 159497 298324 305186
rect 298388 245585 298416 305390
rect 298374 245576 298430 245585
rect 298374 245511 298430 245520
rect 298376 189916 298428 189922
rect 298376 189858 298428 189864
rect 298282 159488 298338 159497
rect 298282 159423 298338 159432
rect 298388 154834 298416 189858
rect 298480 159633 298508 306410
rect 298572 306406 298600 310420
rect 298560 306400 298612 306406
rect 298560 306342 298612 306348
rect 298756 305250 298784 310420
rect 298940 308145 298968 310420
rect 298926 308136 298982 308145
rect 298926 308071 298982 308080
rect 299124 307873 299152 310420
rect 299110 307864 299166 307873
rect 299110 307799 299166 307808
rect 299308 305454 299336 310420
rect 299492 306354 299520 310420
rect 299676 306626 299704 310420
rect 299860 306746 299888 310420
rect 299848 306740 299900 306746
rect 299848 306682 299900 306688
rect 299676 306598 299980 306626
rect 299848 306468 299900 306474
rect 299848 306410 299900 306416
rect 299492 306326 299796 306354
rect 299296 305448 299348 305454
rect 299296 305390 299348 305396
rect 299664 305448 299716 305454
rect 299664 305390 299716 305396
rect 299572 305380 299624 305386
rect 299572 305322 299624 305328
rect 299480 305312 299532 305318
rect 299480 305254 299532 305260
rect 298744 305244 298796 305250
rect 298744 305186 298796 305192
rect 299296 250300 299348 250306
rect 299296 250242 299348 250248
rect 298836 248328 298888 248334
rect 298836 248270 298888 248276
rect 298558 247344 298614 247353
rect 298558 247279 298614 247288
rect 298572 247110 298600 247279
rect 298560 247104 298612 247110
rect 298560 247046 298612 247052
rect 298744 245608 298796 245614
rect 298744 245550 298796 245556
rect 298560 170604 298612 170610
rect 298560 170546 298612 170552
rect 298466 159624 298522 159633
rect 298466 159559 298522 159568
rect 298376 154828 298428 154834
rect 298376 154770 298428 154776
rect 298572 154426 298600 170546
rect 298560 154420 298612 154426
rect 298560 154362 298612 154368
rect 298192 152516 298244 152522
rect 298192 152458 298244 152464
rect 298100 10328 298152 10334
rect 298100 10270 298152 10276
rect 296720 6520 296772 6526
rect 296720 6462 296772 6468
rect 297272 5500 297324 5506
rect 297272 5442 297324 5448
rect 296628 3732 296680 3738
rect 296628 3674 296680 3680
rect 296076 3528 296128 3534
rect 296076 3470 296128 3476
rect 295984 3392 296036 3398
rect 295984 3334 296036 3340
rect 296088 480 296116 3470
rect 297284 480 297312 5442
rect 297364 5228 297416 5234
rect 297364 5170 297416 5176
rect 297376 5030 297404 5170
rect 298468 5092 298520 5098
rect 298468 5034 298520 5040
rect 297364 5024 297416 5030
rect 297364 4966 297416 4972
rect 297456 4072 297508 4078
rect 297456 4014 297508 4020
rect 297468 3602 297496 4014
rect 298100 3800 298152 3806
rect 298100 3742 298152 3748
rect 297456 3596 297508 3602
rect 297456 3538 297508 3544
rect 298112 3330 298140 3742
rect 298100 3324 298152 3330
rect 298100 3266 298152 3272
rect 298480 480 298508 5034
rect 298756 4078 298784 245550
rect 298848 196042 298876 248270
rect 299020 246152 299072 246158
rect 299020 246094 299072 246100
rect 298836 196036 298888 196042
rect 298836 195978 298888 195984
rect 299032 192817 299060 246094
rect 299112 244724 299164 244730
rect 299112 244666 299164 244672
rect 299018 192808 299074 192817
rect 299018 192743 299074 192752
rect 299032 191894 299060 192743
rect 299020 191888 299072 191894
rect 299020 191830 299072 191836
rect 299124 188193 299152 244666
rect 299204 243772 299256 243778
rect 299204 243714 299256 243720
rect 299110 188184 299166 188193
rect 299110 188119 299166 188128
rect 299216 158370 299244 243714
rect 299308 159118 299336 250242
rect 299492 245449 299520 305254
rect 299478 245440 299534 245449
rect 299478 245375 299534 245384
rect 299584 244633 299612 305322
rect 299676 244905 299704 305390
rect 299768 245313 299796 306326
rect 299754 245304 299810 245313
rect 299754 245239 299810 245248
rect 299662 244896 299718 244905
rect 299662 244831 299718 244840
rect 299860 244662 299888 306410
rect 299952 305266 299980 306598
rect 300044 305454 300072 310420
rect 300032 305448 300084 305454
rect 300032 305390 300084 305396
rect 299952 305238 300072 305266
rect 299940 305176 299992 305182
rect 299940 305118 299992 305124
rect 299952 247897 299980 305118
rect 300044 248169 300072 305238
rect 300228 296714 300256 310420
rect 300412 305318 300440 310420
rect 300596 305386 300624 310420
rect 300584 305380 300636 305386
rect 300584 305322 300636 305328
rect 300400 305312 300452 305318
rect 300400 305254 300452 305260
rect 300780 305182 300808 310420
rect 300860 306468 300912 306474
rect 300860 306410 300912 306416
rect 300768 305176 300820 305182
rect 300768 305118 300820 305124
rect 300136 296686 300256 296714
rect 300136 248305 300164 296686
rect 300122 248296 300178 248305
rect 300122 248231 300178 248240
rect 300030 248160 300086 248169
rect 300030 248095 300086 248104
rect 299938 247888 299994 247897
rect 299938 247823 299994 247832
rect 300872 244934 300900 306410
rect 300860 244928 300912 244934
rect 300860 244870 300912 244876
rect 299848 244656 299900 244662
rect 299570 244624 299626 244633
rect 299848 244598 299900 244604
rect 299570 244559 299626 244568
rect 300964 244526 300992 310420
rect 301044 306400 301096 306406
rect 301044 306342 301096 306348
rect 301056 245342 301084 306342
rect 301148 306218 301176 310420
rect 301332 306354 301360 310420
rect 301516 306406 301544 310420
rect 301504 306400 301556 306406
rect 301332 306326 301452 306354
rect 301504 306342 301556 306348
rect 301148 306190 301360 306218
rect 301228 305448 301280 305454
rect 301228 305390 301280 305396
rect 301136 305380 301188 305386
rect 301136 305322 301188 305328
rect 301044 245336 301096 245342
rect 301044 245278 301096 245284
rect 300952 244520 301004 244526
rect 300952 244462 301004 244468
rect 301148 244458 301176 305322
rect 301240 245177 301268 305390
rect 301226 245168 301282 245177
rect 301226 245103 301282 245112
rect 301136 244452 301188 244458
rect 301136 244394 301188 244400
rect 301332 244361 301360 306190
rect 301424 247489 301452 306326
rect 301700 305386 301728 310420
rect 301884 305454 301912 310420
rect 302068 306474 302096 310420
rect 302056 306468 302108 306474
rect 302056 306410 302108 306416
rect 301872 305448 301924 305454
rect 301872 305390 301924 305396
rect 301688 305380 301740 305386
rect 301688 305322 301740 305328
rect 301410 247480 301466 247489
rect 301410 247415 301466 247424
rect 302252 245070 302280 310420
rect 302332 308440 302384 308446
rect 302332 308382 302384 308388
rect 302344 245546 302372 308382
rect 302436 307986 302464 310420
rect 302620 308446 302648 310420
rect 302608 308440 302660 308446
rect 302608 308382 302660 308388
rect 302700 308440 302752 308446
rect 302700 308382 302752 308388
rect 302436 307958 302556 307986
rect 302424 307828 302476 307834
rect 302424 307770 302476 307776
rect 302332 245540 302384 245546
rect 302332 245482 302384 245488
rect 302436 245410 302464 307770
rect 302528 247625 302556 307958
rect 302608 307896 302660 307902
rect 302608 307838 302660 307844
rect 302620 247926 302648 307838
rect 302608 247920 302660 247926
rect 302608 247862 302660 247868
rect 302712 247790 302740 308382
rect 302804 308156 302832 310420
rect 302988 308446 303016 310420
rect 302976 308440 303028 308446
rect 302976 308382 303028 308388
rect 302804 308128 302924 308156
rect 302792 307964 302844 307970
rect 302792 307906 302844 307912
rect 302804 247858 302832 307906
rect 302896 247994 302924 308128
rect 303172 307834 303200 310420
rect 303356 307902 303384 310420
rect 303540 307970 303568 310420
rect 303724 308156 303752 310420
rect 303804 308440 303856 308446
rect 303804 308382 303856 308388
rect 303632 308128 303752 308156
rect 303528 307964 303580 307970
rect 303528 307906 303580 307912
rect 303344 307896 303396 307902
rect 303344 307838 303396 307844
rect 303160 307828 303212 307834
rect 303160 307770 303212 307776
rect 302884 247988 302936 247994
rect 302884 247930 302936 247936
rect 302792 247852 302844 247858
rect 302792 247794 302844 247800
rect 302700 247784 302752 247790
rect 302700 247726 302752 247732
rect 302514 247616 302570 247625
rect 302514 247551 302570 247560
rect 302424 245404 302476 245410
rect 302424 245346 302476 245352
rect 303632 245206 303660 308128
rect 303712 307896 303764 307902
rect 303712 307838 303764 307844
rect 303724 245478 303752 307838
rect 303712 245472 303764 245478
rect 303712 245414 303764 245420
rect 303620 245200 303672 245206
rect 303620 245142 303672 245148
rect 302240 245064 302292 245070
rect 302240 245006 302292 245012
rect 303816 244497 303844 308382
rect 303908 308156 303936 310420
rect 304092 308156 304120 310420
rect 303908 308128 304028 308156
rect 304092 308128 304212 308156
rect 303896 307964 303948 307970
rect 303896 307906 303948 307912
rect 303908 247353 303936 307906
rect 304000 248402 304028 308128
rect 304080 308032 304132 308038
rect 304080 307974 304132 307980
rect 303988 248396 304040 248402
rect 303988 248338 304040 248344
rect 304092 247722 304120 307974
rect 304184 248062 304212 308128
rect 304276 307902 304304 310420
rect 304460 307970 304488 310420
rect 304644 308038 304672 310420
rect 304828 308446 304856 310420
rect 304816 308440 304868 308446
rect 304816 308382 304868 308388
rect 305012 308394 305040 310420
rect 305196 308530 305224 310420
rect 305380 309194 305408 310420
rect 305368 309188 305420 309194
rect 305368 309130 305420 309136
rect 305196 308502 305408 308530
rect 305276 308440 305328 308446
rect 305012 308366 305224 308394
rect 305276 308382 305328 308388
rect 305000 308304 305052 308310
rect 305000 308246 305052 308252
rect 304632 308032 304684 308038
rect 304632 307974 304684 307980
rect 304448 307964 304500 307970
rect 304448 307906 304500 307912
rect 304264 307896 304316 307902
rect 304264 307838 304316 307844
rect 304172 248056 304224 248062
rect 304172 247998 304224 248004
rect 304080 247716 304132 247722
rect 304080 247658 304132 247664
rect 303894 247344 303950 247353
rect 303894 247279 303950 247288
rect 305012 245274 305040 308246
rect 305092 308168 305144 308174
rect 305092 308110 305144 308116
rect 305104 245478 305132 308110
rect 305092 245472 305144 245478
rect 305092 245414 305144 245420
rect 305000 245268 305052 245274
rect 305000 245210 305052 245216
rect 305196 245138 305224 308366
rect 305288 245206 305316 308382
rect 305380 247994 305408 308502
rect 305564 308310 305592 310420
rect 305552 308304 305604 308310
rect 305552 308246 305604 308252
rect 305748 308156 305776 310420
rect 305932 308174 305960 310420
rect 306116 308446 306144 310420
rect 306196 309188 306248 309194
rect 306196 309130 306248 309136
rect 306208 308446 306236 309130
rect 306104 308440 306156 308446
rect 306104 308382 306156 308388
rect 306196 308440 306248 308446
rect 306196 308382 306248 308388
rect 305472 308128 305776 308156
rect 305920 308168 305972 308174
rect 305368 247988 305420 247994
rect 305368 247930 305420 247936
rect 305472 247858 305500 308128
rect 305920 308110 305972 308116
rect 306300 296714 306328 310420
rect 306380 308100 306432 308106
rect 306380 308042 306432 308048
rect 305564 296686 306328 296714
rect 305564 248062 305592 296686
rect 305552 248056 305604 248062
rect 305552 247998 305604 248004
rect 305460 247852 305512 247858
rect 305460 247794 305512 247800
rect 306392 245313 306420 308042
rect 306484 245546 306512 310420
rect 306564 308304 306616 308310
rect 306564 308246 306616 308252
rect 306668 308258 306696 310420
rect 306472 245540 306524 245546
rect 306472 245482 306524 245488
rect 306576 245342 306604 308246
rect 306668 308230 306788 308258
rect 306656 308168 306708 308174
rect 306656 308110 306708 308116
rect 306668 245410 306696 308110
rect 306760 245614 306788 308230
rect 306852 247790 306880 310420
rect 307036 308174 307064 310420
rect 307220 308310 307248 310420
rect 307208 308304 307260 308310
rect 307208 308246 307260 308252
rect 307024 308168 307076 308174
rect 307024 308110 307076 308116
rect 307404 296714 307432 310420
rect 307588 308106 307616 310420
rect 307772 308394 307800 310420
rect 307956 308530 307984 310420
rect 307956 308502 308076 308530
rect 307772 308366 307984 308394
rect 307576 308100 307628 308106
rect 307576 308042 307628 308048
rect 307852 308100 307904 308106
rect 307852 308042 307904 308048
rect 307760 308032 307812 308038
rect 307760 307974 307812 307980
rect 306944 296686 307432 296714
rect 306944 247926 306972 296686
rect 307772 248169 307800 307974
rect 307864 253230 307892 308042
rect 307852 253224 307904 253230
rect 307852 253166 307904 253172
rect 307956 248305 307984 308366
rect 308048 308258 308076 308502
rect 308140 308394 308168 310420
rect 308324 308530 308352 310420
rect 308324 308502 308444 308530
rect 308140 308366 308352 308394
rect 308220 308304 308272 308310
rect 308048 308230 308168 308258
rect 308220 308246 308272 308252
rect 308036 308168 308088 308174
rect 308036 308110 308088 308116
rect 308048 261497 308076 308110
rect 308140 271386 308168 308230
rect 308232 287774 308260 308246
rect 308324 297401 308352 308366
rect 308416 308174 308444 308502
rect 308404 308168 308456 308174
rect 308404 308110 308456 308116
rect 308508 301578 308536 310420
rect 308692 308310 308720 310420
rect 308680 308304 308732 308310
rect 308680 308246 308732 308252
rect 308876 308038 308904 310420
rect 309060 308106 309088 310420
rect 309140 309188 309192 309194
rect 309140 309130 309192 309136
rect 309152 308394 309180 309130
rect 309244 308666 309272 310420
rect 309428 309194 309456 310420
rect 309416 309188 309468 309194
rect 309416 309130 309468 309136
rect 309244 308638 309456 308666
rect 309152 308366 309272 308394
rect 309140 308304 309192 308310
rect 309140 308246 309192 308252
rect 309048 308100 309100 308106
rect 309048 308042 309100 308048
rect 308864 308032 308916 308038
rect 308864 307974 308916 307980
rect 308496 301572 308548 301578
rect 308496 301514 308548 301520
rect 308310 297392 308366 297401
rect 308310 297327 308366 297336
rect 308220 287768 308272 287774
rect 308220 287710 308272 287716
rect 308128 271380 308180 271386
rect 308128 271322 308180 271328
rect 308034 261488 308090 261497
rect 308034 261423 308090 261432
rect 307942 248296 307998 248305
rect 307942 248231 307998 248240
rect 307758 248160 307814 248169
rect 307758 248095 307814 248104
rect 306932 247920 306984 247926
rect 306932 247862 306984 247868
rect 306840 247784 306892 247790
rect 306840 247726 306892 247732
rect 309152 246634 309180 308246
rect 309244 249286 309272 308366
rect 309324 308168 309376 308174
rect 309324 308110 309376 308116
rect 309336 279546 309364 308110
rect 309428 280906 309456 308638
rect 309612 308394 309640 310420
rect 309520 308366 309640 308394
rect 309520 286482 309548 308366
rect 309796 308258 309824 310420
rect 309980 308310 310008 310420
rect 309612 308230 309824 308258
rect 309968 308304 310020 308310
rect 309968 308246 310020 308252
rect 309508 286476 309560 286482
rect 309508 286418 309560 286424
rect 309612 286414 309640 308230
rect 310164 300286 310192 310420
rect 310348 308174 310376 310420
rect 310336 308168 310388 308174
rect 310336 308110 310388 308116
rect 310532 308122 310560 310420
rect 310716 308310 310744 310420
rect 310704 308304 310756 308310
rect 310704 308246 310756 308252
rect 310900 308258 310928 310420
rect 310900 308230 311020 308258
rect 310532 308094 310928 308122
rect 310612 308032 310664 308038
rect 310612 307974 310664 307980
rect 310520 307828 310572 307834
rect 310520 307770 310572 307776
rect 310152 300280 310204 300286
rect 310152 300222 310204 300228
rect 309600 286408 309652 286414
rect 309600 286350 309652 286356
rect 309416 280900 309468 280906
rect 309416 280842 309468 280848
rect 309324 279540 309376 279546
rect 309324 279482 309376 279488
rect 310532 250578 310560 307770
rect 310624 250646 310652 307974
rect 310704 307964 310756 307970
rect 310704 307906 310756 307912
rect 310716 278118 310744 307906
rect 310796 307896 310848 307902
rect 310796 307838 310848 307844
rect 310808 282266 310836 307838
rect 310900 282334 310928 308094
rect 310992 294846 311020 308230
rect 311084 308038 311112 310420
rect 311072 308032 311124 308038
rect 311072 307974 311124 307980
rect 311268 303249 311296 310420
rect 311452 307970 311480 310420
rect 311440 307964 311492 307970
rect 311440 307906 311492 307912
rect 311636 307834 311664 310420
rect 311716 308304 311768 308310
rect 311716 308246 311768 308252
rect 311728 308038 311756 308246
rect 311716 308032 311768 308038
rect 311716 307974 311768 307980
rect 311820 307902 311848 310420
rect 311808 307896 311860 307902
rect 311808 307838 311860 307844
rect 311624 307828 311676 307834
rect 311624 307770 311676 307776
rect 311900 306400 311952 306406
rect 311900 306342 311952 306348
rect 311254 303240 311310 303249
rect 311254 303175 311310 303184
rect 310980 294840 311032 294846
rect 310980 294782 311032 294788
rect 310888 282328 310940 282334
rect 310888 282270 310940 282276
rect 310796 282260 310848 282266
rect 310796 282202 310848 282208
rect 310704 278112 310756 278118
rect 310704 278054 310756 278060
rect 310612 250640 310664 250646
rect 310612 250582 310664 250588
rect 310520 250572 310572 250578
rect 310520 250514 310572 250520
rect 309232 249280 309284 249286
rect 309232 249222 309284 249228
rect 309140 246628 309192 246634
rect 309140 246570 309192 246576
rect 306748 245608 306800 245614
rect 306748 245550 306800 245556
rect 306656 245404 306708 245410
rect 306656 245346 306708 245352
rect 306564 245336 306616 245342
rect 306378 245304 306434 245313
rect 306564 245278 306616 245284
rect 306378 245239 306434 245248
rect 305276 245200 305328 245206
rect 305276 245142 305328 245148
rect 305184 245132 305236 245138
rect 305184 245074 305236 245080
rect 311912 245070 311940 306342
rect 312004 303906 312032 310420
rect 312188 306406 312216 310420
rect 312176 306400 312228 306406
rect 312176 306342 312228 306348
rect 312004 303878 312308 303906
rect 312176 303816 312228 303822
rect 312176 303758 312228 303764
rect 311992 303748 312044 303754
rect 311992 303690 312044 303696
rect 312004 260370 312032 303690
rect 312084 303680 312136 303686
rect 312084 303622 312136 303628
rect 312096 273970 312124 303622
rect 312188 275398 312216 303758
rect 312280 276758 312308 303878
rect 312372 298858 312400 310420
rect 312452 308032 312504 308038
rect 312452 307974 312504 307980
rect 312464 302234 312492 307974
rect 312556 303822 312584 310420
rect 312544 303816 312596 303822
rect 312544 303758 312596 303764
rect 312740 303754 312768 310420
rect 312924 307834 312952 310420
rect 312912 307828 312964 307834
rect 312912 307770 312964 307776
rect 312728 303748 312780 303754
rect 312728 303690 312780 303696
rect 313108 303686 313136 310420
rect 313096 303680 313148 303686
rect 313096 303622 313148 303628
rect 312464 302206 312584 302234
rect 312360 298852 312412 298858
rect 312360 298794 312412 298800
rect 312556 285122 312584 302206
rect 312544 285116 312596 285122
rect 312544 285058 312596 285064
rect 312268 276752 312320 276758
rect 312268 276694 312320 276700
rect 312176 275392 312228 275398
rect 312176 275334 312228 275340
rect 312084 273964 312136 273970
rect 312084 273906 312136 273912
rect 311992 260364 312044 260370
rect 311992 260306 312044 260312
rect 313292 258942 313320 310420
rect 313372 306400 313424 306406
rect 313372 306342 313424 306348
rect 313384 268734 313412 306342
rect 313476 304722 313504 310420
rect 313660 305386 313688 310420
rect 313844 306354 313872 310420
rect 314028 306406 314056 310420
rect 313752 306326 313872 306354
rect 314016 306400 314068 306406
rect 314016 306342 314068 306348
rect 313648 305380 313700 305386
rect 313648 305322 313700 305328
rect 313476 304694 313688 304722
rect 313556 304632 313608 304638
rect 313556 304574 313608 304580
rect 313464 304564 313516 304570
rect 313464 304506 313516 304512
rect 313372 268728 313424 268734
rect 313372 268670 313424 268676
rect 313476 268666 313504 304506
rect 313568 271318 313596 304574
rect 313660 283694 313688 304694
rect 313648 283688 313700 283694
rect 313648 283630 313700 283636
rect 313752 283626 313780 306326
rect 313832 305380 313884 305386
rect 313832 305322 313884 305328
rect 313844 285054 313872 305322
rect 314212 304638 314240 310420
rect 314200 304632 314252 304638
rect 314200 304574 314252 304580
rect 314396 304570 314424 310420
rect 314384 304564 314436 304570
rect 314384 304506 314436 304512
rect 314580 296714 314608 310420
rect 314764 307154 314792 310420
rect 314752 307148 314804 307154
rect 314752 307090 314804 307096
rect 314752 306536 314804 306542
rect 314752 306478 314804 306484
rect 314660 306400 314712 306406
rect 314660 306342 314712 306348
rect 313936 296686 314608 296714
rect 313936 291922 313964 296686
rect 313924 291916 313976 291922
rect 313924 291858 313976 291864
rect 313832 285048 313884 285054
rect 313832 284990 313884 284996
rect 313740 283620 313792 283626
rect 313740 283562 313792 283568
rect 313556 271312 313608 271318
rect 313556 271254 313608 271260
rect 313464 268660 313516 268666
rect 313464 268602 313516 268608
rect 313280 258936 313332 258942
rect 313280 258878 313332 258884
rect 314672 249218 314700 306342
rect 314764 267170 314792 306478
rect 314844 306468 314896 306474
rect 314844 306410 314896 306416
rect 314856 268598 314884 306410
rect 314948 270026 314976 310420
rect 315132 306406 315160 310420
rect 315316 308122 315344 310420
rect 315316 308094 315436 308122
rect 315304 307828 315356 307834
rect 315304 307770 315356 307776
rect 315120 306400 315172 306406
rect 315120 306342 315172 306348
rect 314936 270020 314988 270026
rect 314936 269962 314988 269968
rect 314844 268592 314896 268598
rect 314844 268534 314896 268540
rect 314752 267164 314804 267170
rect 314752 267106 314804 267112
rect 315316 252006 315344 307770
rect 315408 305969 315436 308094
rect 315500 306474 315528 310420
rect 315684 306542 315712 310420
rect 315672 306536 315724 306542
rect 315672 306478 315724 306484
rect 315488 306468 315540 306474
rect 315488 306410 315540 306416
rect 315394 305960 315450 305969
rect 315394 305895 315450 305904
rect 315868 304366 315896 310420
rect 316052 306354 316080 310420
rect 316236 307086 316264 310420
rect 316224 307080 316276 307086
rect 316224 307022 316276 307028
rect 316224 306468 316276 306474
rect 316224 306410 316276 306416
rect 316052 306326 316172 306354
rect 316040 305380 316092 305386
rect 316040 305322 316092 305328
rect 315856 304360 315908 304366
rect 315856 304302 315908 304308
rect 315304 252000 315356 252006
rect 315304 251942 315356 251948
rect 314660 249212 314712 249218
rect 314660 249154 314712 249160
rect 316052 246566 316080 305322
rect 316144 258874 316172 306326
rect 316132 258868 316184 258874
rect 316132 258810 316184 258816
rect 316236 258806 316264 306410
rect 316420 305386 316448 310420
rect 316604 306474 316632 310420
rect 316592 306468 316644 306474
rect 316592 306410 316644 306416
rect 316788 306354 316816 310420
rect 316868 307964 316920 307970
rect 316868 307906 316920 307912
rect 316512 306326 316816 306354
rect 316408 305380 316460 305386
rect 316408 305322 316460 305328
rect 316316 305312 316368 305318
rect 316316 305254 316368 305260
rect 316328 260302 316356 305254
rect 316408 305244 316460 305250
rect 316408 305186 316460 305192
rect 316420 265742 316448 305186
rect 316512 267102 316540 306326
rect 316880 302234 316908 307906
rect 316972 305833 317000 310420
rect 316958 305824 317014 305833
rect 316958 305759 317014 305768
rect 317156 305318 317184 310420
rect 317144 305312 317196 305318
rect 317144 305254 317196 305260
rect 317340 305250 317368 310420
rect 317524 306542 317552 310420
rect 317512 306536 317564 306542
rect 317512 306478 317564 306484
rect 317512 306400 317564 306406
rect 317708 306354 317736 310420
rect 317512 306342 317564 306348
rect 317328 305244 317380 305250
rect 317328 305186 317380 305192
rect 317420 304428 317472 304434
rect 317420 304370 317472 304376
rect 316788 302206 316908 302234
rect 316500 267096 316552 267102
rect 316500 267038 316552 267044
rect 316408 265736 316460 265742
rect 316408 265678 316460 265684
rect 316316 260296 316368 260302
rect 316316 260238 316368 260244
rect 316224 258800 316276 258806
rect 316224 258742 316276 258748
rect 316040 246560 316092 246566
rect 316040 246502 316092 246508
rect 311900 245064 311952 245070
rect 311900 245006 311952 245012
rect 303802 244488 303858 244497
rect 303802 244423 303858 244432
rect 301318 244352 301374 244361
rect 301318 244287 301374 244296
rect 316788 243846 316816 302206
rect 317432 264382 317460 304370
rect 317524 265674 317552 306342
rect 317616 306326 317736 306354
rect 317616 267034 317644 306326
rect 317892 306218 317920 310420
rect 317972 306536 318024 306542
rect 317972 306478 318024 306484
rect 317708 306190 317920 306218
rect 317708 279478 317736 306190
rect 317788 305380 317840 305386
rect 317788 305322 317840 305328
rect 317800 300218 317828 305322
rect 317984 303113 318012 306478
rect 317970 303104 318026 303113
rect 317970 303039 318026 303048
rect 318076 302234 318104 310420
rect 318260 306406 318288 310420
rect 318248 306400 318300 306406
rect 318248 306342 318300 306348
rect 318444 304434 318472 310420
rect 318628 305386 318656 310420
rect 318616 305380 318668 305386
rect 318616 305322 318668 305328
rect 318812 305318 318840 310420
rect 318892 306400 318944 306406
rect 318892 306342 318944 306348
rect 318800 305312 318852 305318
rect 318800 305254 318852 305260
rect 318800 305176 318852 305182
rect 318800 305118 318852 305124
rect 318432 304428 318484 304434
rect 318432 304370 318484 304376
rect 317892 302206 318104 302234
rect 317892 301510 317920 302206
rect 317880 301504 317932 301510
rect 317880 301446 317932 301452
rect 317788 300212 317840 300218
rect 317788 300154 317840 300160
rect 317696 279472 317748 279478
rect 317696 279414 317748 279420
rect 317604 267028 317656 267034
rect 317604 266970 317656 266976
rect 317512 265668 317564 265674
rect 317512 265610 317564 265616
rect 317420 264376 317472 264382
rect 317420 264318 317472 264324
rect 318812 250510 318840 305118
rect 318904 263158 318932 306342
rect 318996 305386 319024 310420
rect 319076 306876 319128 306882
rect 319076 306818 319128 306824
rect 318984 305380 319036 305386
rect 318984 305322 319036 305328
rect 318984 305244 319036 305250
rect 318984 305186 319036 305192
rect 318996 264314 319024 305186
rect 319088 280838 319116 306818
rect 319180 306388 319208 310420
rect 319364 306882 319392 310420
rect 319352 306876 319404 306882
rect 319352 306818 319404 306824
rect 319548 306406 319576 310420
rect 319536 306400 319588 306406
rect 319180 306360 319392 306388
rect 319260 305380 319312 305386
rect 319260 305322 319312 305328
rect 319168 305312 319220 305318
rect 319168 305254 319220 305260
rect 319180 282198 319208 305254
rect 319272 294778 319300 305322
rect 319364 304298 319392 306360
rect 319536 306342 319588 306348
rect 319352 304292 319404 304298
rect 319352 304234 319404 304240
rect 319732 302234 319760 310420
rect 319916 305250 319944 310420
rect 319904 305244 319956 305250
rect 319904 305186 319956 305192
rect 320100 305182 320128 310420
rect 320284 306474 320312 310420
rect 320272 306468 320324 306474
rect 320272 306410 320324 306416
rect 320180 306400 320232 306406
rect 320468 306354 320496 310420
rect 320180 306342 320232 306348
rect 320088 305176 320140 305182
rect 320088 305118 320140 305124
rect 319364 302206 319760 302234
rect 319364 298790 319392 302206
rect 319352 298784 319404 298790
rect 319352 298726 319404 298732
rect 319260 294772 319312 294778
rect 319260 294714 319312 294720
rect 319168 282192 319220 282198
rect 319168 282134 319220 282140
rect 319076 280832 319128 280838
rect 319076 280774 319128 280780
rect 318984 264308 319036 264314
rect 318984 264250 319036 264256
rect 318892 263152 318944 263158
rect 318892 263094 318944 263100
rect 320192 261730 320220 306342
rect 320284 306326 320496 306354
rect 320284 263090 320312 306326
rect 320652 306218 320680 310420
rect 320732 306468 320784 306474
rect 320732 306410 320784 306416
rect 320468 306190 320680 306218
rect 320364 305312 320416 305318
rect 320364 305254 320416 305260
rect 320376 276690 320404 305254
rect 320468 278050 320496 306190
rect 320548 305380 320600 305386
rect 320548 305322 320600 305328
rect 320560 296070 320588 305322
rect 320744 302977 320772 306410
rect 320730 302968 320786 302977
rect 320730 302903 320786 302912
rect 320836 302234 320864 310420
rect 321020 306406 321048 310420
rect 321008 306400 321060 306406
rect 321008 306342 321060 306348
rect 321204 305318 321232 310420
rect 321388 305386 321416 310420
rect 321572 308530 321600 310420
rect 321480 308502 321600 308530
rect 321480 308242 321508 308502
rect 321468 308236 321520 308242
rect 321468 308178 321520 308184
rect 321756 306474 321784 310420
rect 321836 308236 321888 308242
rect 321836 308178 321888 308184
rect 321744 306468 321796 306474
rect 321744 306410 321796 306416
rect 321560 306400 321612 306406
rect 321560 306342 321612 306348
rect 321376 305380 321428 305386
rect 321376 305322 321428 305328
rect 321192 305312 321244 305318
rect 321192 305254 321244 305260
rect 320652 302206 320864 302234
rect 320652 297430 320680 302206
rect 320640 297424 320692 297430
rect 320640 297366 320692 297372
rect 320548 296064 320600 296070
rect 320548 296006 320600 296012
rect 320456 278044 320508 278050
rect 320456 277986 320508 277992
rect 320364 276684 320416 276690
rect 320364 276626 320416 276632
rect 320272 263084 320324 263090
rect 320272 263026 320324 263032
rect 320180 261724 320232 261730
rect 320180 261666 320232 261672
rect 318800 250504 318852 250510
rect 318800 250446 318852 250452
rect 321572 245002 321600 306342
rect 321848 306218 321876 308178
rect 321940 306406 321968 310420
rect 321928 306400 321980 306406
rect 322124 306354 322152 310420
rect 322204 306468 322256 306474
rect 322204 306410 322256 306416
rect 321928 306342 321980 306348
rect 322032 306326 322152 306354
rect 321848 306190 321968 306218
rect 321836 305380 321888 305386
rect 321836 305322 321888 305328
rect 321652 305312 321704 305318
rect 321652 305254 321704 305260
rect 321664 248033 321692 305254
rect 321744 305244 321796 305250
rect 321744 305186 321796 305192
rect 321756 251870 321784 305186
rect 321848 251938 321876 305322
rect 321940 257378 321968 306190
rect 322032 260234 322060 306326
rect 322112 305176 322164 305182
rect 322112 305118 322164 305124
rect 322124 261662 322152 305118
rect 322216 268530 322244 306410
rect 322308 305386 322336 310420
rect 322296 305380 322348 305386
rect 322296 305322 322348 305328
rect 322492 305318 322520 310420
rect 322480 305312 322532 305318
rect 322480 305254 322532 305260
rect 322676 305182 322704 310420
rect 322860 305250 322888 310420
rect 323044 306490 323072 310420
rect 322952 306462 323072 306490
rect 322952 305318 322980 306462
rect 323228 306354 323256 310420
rect 323412 306490 323440 310420
rect 323044 306326 323256 306354
rect 323320 306462 323440 306490
rect 322940 305312 322992 305318
rect 322940 305254 322992 305260
rect 322848 305244 322900 305250
rect 322848 305186 322900 305192
rect 322664 305176 322716 305182
rect 322664 305118 322716 305124
rect 322940 305176 322992 305182
rect 322940 305118 322992 305124
rect 322204 268524 322256 268530
rect 322204 268466 322256 268472
rect 322112 261656 322164 261662
rect 322112 261598 322164 261604
rect 322020 260228 322072 260234
rect 322020 260170 322072 260176
rect 321928 257372 321980 257378
rect 321928 257314 321980 257320
rect 321836 251932 321888 251938
rect 321836 251874 321888 251880
rect 321744 251864 321796 251870
rect 321744 251806 321796 251812
rect 321650 248024 321706 248033
rect 321650 247959 321706 247968
rect 322952 246498 322980 305118
rect 323044 247897 323072 306326
rect 323320 306218 323348 306462
rect 323596 306354 323624 310420
rect 323136 306190 323348 306218
rect 323412 306326 323624 306354
rect 323136 261594 323164 306190
rect 323308 305380 323360 305386
rect 323308 305322 323360 305328
rect 323216 305244 323268 305250
rect 323216 305186 323268 305192
rect 323228 275330 323256 305186
rect 323320 291854 323348 305322
rect 323412 293350 323440 306326
rect 323492 305312 323544 305318
rect 323492 305254 323544 305260
rect 323504 294710 323532 305254
rect 323780 305182 323808 310420
rect 323964 305250 323992 310420
rect 324148 305386 324176 310420
rect 324332 306354 324360 310420
rect 324516 306474 324544 310420
rect 324700 306626 324728 310420
rect 324608 306598 324728 306626
rect 324504 306468 324556 306474
rect 324504 306410 324556 306416
rect 324332 306326 324544 306354
rect 324410 305688 324466 305697
rect 324410 305623 324466 305632
rect 324136 305380 324188 305386
rect 324136 305322 324188 305328
rect 324320 305380 324372 305386
rect 324320 305322 324372 305328
rect 323952 305244 324004 305250
rect 323952 305186 324004 305192
rect 323768 305176 323820 305182
rect 323768 305118 323820 305124
rect 323492 294704 323544 294710
rect 323492 294646 323544 294652
rect 323400 293344 323452 293350
rect 323400 293286 323452 293292
rect 323308 291848 323360 291854
rect 323308 291790 323360 291796
rect 323216 275324 323268 275330
rect 323216 275266 323268 275272
rect 323124 261588 323176 261594
rect 323124 261530 323176 261536
rect 323030 247888 323086 247897
rect 323030 247823 323086 247832
rect 322940 246492 322992 246498
rect 322940 246434 322992 246440
rect 324332 246430 324360 305322
rect 324424 247761 324452 305623
rect 324516 261526 324544 306326
rect 324608 305386 324636 306598
rect 324884 306490 324912 310420
rect 324700 306462 324912 306490
rect 324596 305380 324648 305386
rect 324596 305322 324648 305328
rect 324596 305244 324648 305250
rect 324596 305186 324648 305192
rect 324608 262954 324636 305186
rect 324700 263022 324728 306462
rect 325068 306354 325096 310420
rect 325148 306468 325200 306474
rect 325148 306410 325200 306416
rect 324792 306326 325096 306354
rect 324792 268462 324820 306326
rect 324872 305380 324924 305386
rect 324872 305322 324924 305328
rect 324780 268456 324832 268462
rect 324780 268398 324832 268404
rect 324884 268394 324912 305322
rect 325160 296714 325188 306410
rect 325252 305697 325280 310420
rect 325238 305688 325294 305697
rect 325238 305623 325294 305632
rect 325436 305250 325464 310420
rect 325620 305386 325648 310420
rect 325804 306354 325832 310420
rect 325884 306468 325936 306474
rect 325884 306410 325936 306416
rect 325712 306326 325832 306354
rect 325608 305380 325660 305386
rect 325608 305322 325660 305328
rect 325424 305244 325476 305250
rect 325424 305186 325476 305192
rect 324976 296686 325188 296714
rect 324976 294642 325004 296686
rect 324964 294636 325016 294642
rect 324964 294578 325016 294584
rect 324872 268388 324924 268394
rect 324872 268330 324924 268336
rect 324688 263016 324740 263022
rect 324688 262958 324740 262964
rect 324596 262948 324648 262954
rect 324596 262890 324648 262896
rect 324504 261520 324556 261526
rect 324504 261462 324556 261468
rect 324410 247752 324466 247761
rect 324410 247687 324466 247696
rect 325712 247625 325740 306326
rect 325792 305312 325844 305318
rect 325792 305254 325844 305260
rect 325804 249082 325832 305254
rect 325896 249150 325924 306410
rect 325988 262886 326016 310420
rect 326068 306400 326120 306406
rect 326068 306342 326120 306348
rect 326172 306354 326200 310420
rect 326356 306474 326384 310420
rect 326344 306468 326396 306474
rect 326344 306410 326396 306416
rect 326540 306406 326568 310420
rect 326528 306400 326580 306406
rect 326080 264246 326108 306342
rect 326172 306326 326292 306354
rect 326528 306342 326580 306348
rect 326160 305380 326212 305386
rect 326160 305322 326212 305328
rect 326172 269958 326200 305322
rect 326264 286346 326292 306326
rect 326724 305386 326752 310420
rect 326712 305380 326764 305386
rect 326712 305322 326764 305328
rect 326908 305318 326936 310420
rect 327092 305386 327120 310420
rect 327172 306400 327224 306406
rect 327172 306342 327224 306348
rect 327276 306354 327304 310420
rect 327460 306474 327488 310420
rect 327448 306468 327500 306474
rect 327448 306410 327500 306416
rect 327644 306354 327672 310420
rect 327828 306406 327856 310420
rect 327080 305380 327132 305386
rect 327080 305322 327132 305328
rect 326896 305312 326948 305318
rect 326896 305254 326948 305260
rect 327080 305244 327132 305250
rect 327080 305186 327132 305192
rect 326252 286340 326304 286346
rect 326252 286282 326304 286288
rect 326160 269952 326212 269958
rect 326160 269894 326212 269900
rect 326068 264240 326120 264246
rect 326068 264182 326120 264188
rect 325976 262880 326028 262886
rect 325976 262822 326028 262828
rect 325884 249144 325936 249150
rect 325884 249086 325936 249092
rect 325792 249076 325844 249082
rect 325792 249018 325844 249024
rect 325698 247616 325754 247625
rect 325698 247551 325754 247560
rect 324320 246424 324372 246430
rect 324320 246366 324372 246372
rect 327092 245177 327120 305186
rect 327184 246362 327212 306342
rect 327276 306326 327396 306354
rect 327264 305312 327316 305318
rect 327264 305254 327316 305260
rect 327276 269890 327304 305254
rect 327368 271250 327396 306326
rect 327460 306326 327672 306354
rect 327816 306400 327868 306406
rect 327816 306342 327868 306348
rect 327460 284986 327488 306326
rect 328012 306218 328040 310420
rect 328092 306468 328144 306474
rect 328092 306410 328144 306416
rect 327552 306190 328040 306218
rect 327552 290494 327580 306190
rect 327632 305380 327684 305386
rect 327632 305322 327684 305328
rect 327644 300150 327672 305322
rect 328104 302841 328132 306410
rect 328196 305250 328224 310420
rect 328380 305318 328408 310420
rect 328460 306536 328512 306542
rect 328460 306478 328512 306484
rect 328368 305312 328420 305318
rect 328368 305254 328420 305260
rect 328184 305244 328236 305250
rect 328184 305186 328236 305192
rect 328090 302832 328146 302841
rect 328090 302767 328146 302776
rect 327632 300144 327684 300150
rect 327632 300086 327684 300092
rect 327540 290488 327592 290494
rect 327540 290430 327592 290436
rect 327448 284980 327500 284986
rect 327448 284922 327500 284928
rect 327356 271244 327408 271250
rect 327356 271186 327408 271192
rect 327264 269884 327316 269890
rect 327264 269826 327316 269832
rect 327172 246356 327224 246362
rect 327172 246298 327224 246304
rect 327078 245168 327134 245177
rect 327078 245103 327134 245112
rect 328472 245041 328500 306478
rect 328564 306474 328592 310420
rect 328552 306468 328604 306474
rect 328552 306410 328604 306416
rect 328748 306354 328776 310420
rect 328656 306326 328776 306354
rect 328828 306400 328880 306406
rect 328828 306342 328880 306348
rect 328552 305312 328604 305318
rect 328552 305254 328604 305260
rect 328564 269822 328592 305254
rect 328656 271182 328684 306326
rect 328736 305380 328788 305386
rect 328736 305322 328788 305328
rect 328748 287706 328776 305322
rect 328840 289134 328868 306342
rect 328932 293282 328960 310420
rect 329012 306468 329064 306474
rect 329012 306410 329064 306416
rect 329024 296002 329052 306410
rect 329116 306406 329144 310420
rect 329104 306400 329156 306406
rect 329104 306342 329156 306348
rect 329300 305318 329328 310420
rect 329380 306604 329432 306610
rect 329380 306546 329432 306552
rect 329392 306270 329420 306546
rect 329484 306542 329512 310420
rect 329472 306536 329524 306542
rect 329472 306478 329524 306484
rect 329380 306264 329432 306270
rect 329380 306206 329432 306212
rect 329668 305386 329696 310420
rect 329656 305380 329708 305386
rect 329656 305322 329708 305328
rect 329288 305312 329340 305318
rect 329288 305254 329340 305260
rect 329852 302234 329880 310420
rect 329852 302206 329972 302234
rect 329012 295996 329064 296002
rect 329012 295938 329064 295944
rect 328920 293276 328972 293282
rect 328920 293218 328972 293224
rect 328828 289128 328880 289134
rect 328828 289070 328880 289076
rect 328736 287700 328788 287706
rect 328736 287642 328788 287648
rect 328644 271176 328696 271182
rect 328644 271118 328696 271124
rect 328552 269816 328604 269822
rect 328552 269758 328604 269764
rect 328458 245032 328514 245041
rect 321560 244996 321612 245002
rect 328458 244967 328514 244976
rect 321560 244938 321612 244944
rect 329944 244934 329972 302206
rect 329932 244928 329984 244934
rect 330036 244905 330064 310420
rect 330220 306354 330248 310420
rect 330128 306326 330248 306354
rect 330128 256154 330156 306326
rect 330404 305561 330432 310420
rect 330390 305552 330446 305561
rect 330390 305487 330446 305496
rect 330588 302234 330616 310420
rect 330772 303618 330800 310420
rect 330956 308378 330984 310420
rect 330944 308372 330996 308378
rect 330944 308314 330996 308320
rect 331140 307902 331168 310420
rect 331324 308281 331352 310420
rect 331310 308272 331366 308281
rect 331310 308207 331366 308216
rect 331128 307896 331180 307902
rect 331128 307838 331180 307844
rect 331508 306490 331536 310420
rect 331416 306462 331536 306490
rect 330760 303612 330812 303618
rect 330760 303554 330812 303560
rect 331416 302734 331444 306462
rect 331496 306400 331548 306406
rect 331496 306342 331548 306348
rect 331404 302728 331456 302734
rect 331404 302670 331456 302676
rect 330220 302206 330616 302234
rect 330116 256148 330168 256154
rect 330116 256090 330168 256096
rect 329932 244870 329984 244876
rect 330022 244896 330078 244905
rect 330022 244831 330078 244840
rect 330220 244594 330248 302206
rect 331508 300558 331536 306342
rect 331692 302802 331720 310420
rect 331876 309058 331904 310420
rect 331864 309052 331916 309058
rect 331864 308994 331916 309000
rect 331956 309052 332008 309058
rect 331956 308994 332008 309000
rect 331680 302796 331732 302802
rect 331680 302738 331732 302744
rect 331968 302234 331996 308994
rect 332060 305454 332088 310420
rect 332244 306241 332272 310420
rect 332428 306406 332456 310420
rect 332508 308372 332560 308378
rect 332508 308314 332560 308320
rect 332416 306400 332468 306406
rect 332416 306342 332468 306348
rect 332230 306232 332286 306241
rect 332230 306167 332286 306176
rect 332232 306128 332284 306134
rect 332284 306076 332456 306082
rect 332232 306070 332456 306076
rect 332244 306054 332456 306070
rect 332428 305590 332456 306054
rect 332416 305584 332468 305590
rect 332416 305526 332468 305532
rect 332048 305448 332100 305454
rect 332048 305390 332100 305396
rect 332520 302234 332548 308314
rect 332612 302870 332640 310420
rect 332692 306468 332744 306474
rect 332692 306410 332744 306416
rect 332600 302864 332652 302870
rect 332600 302806 332652 302812
rect 331876 302206 331996 302234
rect 332336 302206 332548 302234
rect 331496 300552 331548 300558
rect 331496 300494 331548 300500
rect 331876 246974 331904 302206
rect 332336 296714 332364 302206
rect 331968 296686 332364 296714
rect 331968 250850 331996 296686
rect 332704 256086 332732 306410
rect 332796 302234 332824 310420
rect 332980 306610 333008 310420
rect 332968 306604 333020 306610
rect 332968 306546 333020 306552
rect 333164 303521 333192 310420
rect 333150 303512 333206 303521
rect 333150 303447 333206 303456
rect 333348 302234 333376 310420
rect 332796 302206 333008 302234
rect 332692 256080 332744 256086
rect 332692 256022 332744 256028
rect 331956 250844 332008 250850
rect 331956 250786 332008 250792
rect 331864 246968 331916 246974
rect 331864 246910 331916 246916
rect 332980 244730 333008 302206
rect 333164 302206 333376 302234
rect 333164 300626 333192 302206
rect 333532 300694 333560 310420
rect 333716 306474 333744 310420
rect 333704 306468 333756 306474
rect 333704 306410 333756 306416
rect 333900 305386 333928 310420
rect 334084 306490 334112 310420
rect 333992 306462 334112 306490
rect 333888 305380 333940 305386
rect 333888 305322 333940 305328
rect 333992 303385 334020 306462
rect 334268 306354 334296 310420
rect 334348 306468 334400 306474
rect 334348 306410 334400 306416
rect 334084 306326 334296 306354
rect 333978 303376 334034 303385
rect 333978 303311 334034 303320
rect 333520 300688 333572 300694
rect 333520 300630 333572 300636
rect 333152 300620 333204 300626
rect 333152 300562 333204 300568
rect 334084 251190 334112 306326
rect 334164 306264 334216 306270
rect 334164 306206 334216 306212
rect 334072 251184 334124 251190
rect 334072 251126 334124 251132
rect 334176 250374 334204 306206
rect 334164 250368 334216 250374
rect 334164 250310 334216 250316
rect 334360 247518 334388 306410
rect 334452 306354 334480 310420
rect 334636 306474 334664 310420
rect 334624 306468 334676 306474
rect 334624 306410 334676 306416
rect 334452 306326 334756 306354
rect 334820 306338 334848 310420
rect 334728 300762 334756 306326
rect 334808 306332 334860 306338
rect 334808 306274 334860 306280
rect 335004 303482 335032 310420
rect 335188 306270 335216 310420
rect 335372 306270 335400 310420
rect 335176 306264 335228 306270
rect 335176 306206 335228 306212
rect 335360 306264 335412 306270
rect 335360 306206 335412 306212
rect 335556 306134 335584 310420
rect 335740 306490 335768 310420
rect 335820 309120 335872 309126
rect 335820 309062 335872 309068
rect 335832 308242 335860 309062
rect 335820 308236 335872 308242
rect 335820 308178 335872 308184
rect 335648 306462 335768 306490
rect 335544 306128 335596 306134
rect 335544 306070 335596 306076
rect 335648 304042 335676 306462
rect 335924 306354 335952 310420
rect 336004 309120 336056 309126
rect 336004 309062 336056 309068
rect 336016 308854 336044 309062
rect 336004 308848 336056 308854
rect 336004 308790 336056 308796
rect 336004 308508 336056 308514
rect 336004 308450 336056 308456
rect 336016 307834 336044 308450
rect 336004 307828 336056 307834
rect 336004 307770 336056 307776
rect 335556 304014 335676 304042
rect 335740 306326 335952 306354
rect 334992 303476 335044 303482
rect 334992 303418 335044 303424
rect 335556 303414 335584 304014
rect 335636 303884 335688 303890
rect 335636 303826 335688 303832
rect 335544 303408 335596 303414
rect 335544 303350 335596 303356
rect 334716 300756 334768 300762
rect 334716 300698 334768 300704
rect 334348 247512 334400 247518
rect 334348 247454 334400 247460
rect 335648 247450 335676 303826
rect 335636 247444 335688 247450
rect 335636 247386 335688 247392
rect 332968 244724 333020 244730
rect 332968 244666 333020 244672
rect 330208 244588 330260 244594
rect 330208 244530 330260 244536
rect 316776 243840 316828 243846
rect 316776 243782 316828 243788
rect 335740 243710 335768 306326
rect 335820 306264 335872 306270
rect 335820 306206 335872 306212
rect 335832 246158 335860 306206
rect 336108 296714 336136 310420
rect 336292 305454 336320 310420
rect 336280 305448 336332 305454
rect 336280 305390 336332 305396
rect 336476 303346 336504 310420
rect 336660 303890 336688 310420
rect 336844 306354 336872 310420
rect 337028 306490 337056 310420
rect 337212 306626 337240 310420
rect 337212 306598 337332 306626
rect 337028 306462 337240 306490
rect 336844 306326 337148 306354
rect 336924 306264 336976 306270
rect 336924 306206 336976 306212
rect 336648 303884 336700 303890
rect 336648 303826 336700 303832
rect 336464 303340 336516 303346
rect 336464 303282 336516 303288
rect 336016 296686 336136 296714
rect 336016 246226 336044 296686
rect 336936 256018 336964 306206
rect 336924 256012 336976 256018
rect 336924 255954 336976 255960
rect 336004 246220 336056 246226
rect 336004 246162 336056 246168
rect 335820 246152 335872 246158
rect 335820 246094 335872 246100
rect 337120 244798 337148 306326
rect 337212 305590 337240 306462
rect 337200 305584 337252 305590
rect 337200 305526 337252 305532
rect 337304 303278 337332 306598
rect 337292 303272 337344 303278
rect 337292 303214 337344 303220
rect 337396 302234 337424 310420
rect 337580 306270 337608 310420
rect 337568 306264 337620 306270
rect 337568 306206 337620 306212
rect 337764 303550 337792 310420
rect 337752 303544 337804 303550
rect 337752 303486 337804 303492
rect 337948 303210 337976 310420
rect 337936 303204 337988 303210
rect 337936 303146 337988 303152
rect 338132 302394 338160 310420
rect 338316 306354 338344 310420
rect 338500 306490 338528 310420
rect 338500 306462 338620 306490
rect 338316 306326 338528 306354
rect 338304 306264 338356 306270
rect 338304 306206 338356 306212
rect 338120 302388 338172 302394
rect 338120 302330 338172 302336
rect 337212 302206 337424 302234
rect 337212 248266 337240 302206
rect 338316 250986 338344 306206
rect 338396 303340 338448 303346
rect 338396 303282 338448 303288
rect 338304 250980 338356 250986
rect 338304 250922 338356 250928
rect 338408 250918 338436 303282
rect 338396 250912 338448 250918
rect 338396 250854 338448 250860
rect 337200 248260 337252 248266
rect 337200 248202 337252 248208
rect 337108 244792 337160 244798
rect 337108 244734 337160 244740
rect 338500 243778 338528 306326
rect 338592 303074 338620 306462
rect 338684 303346 338712 310420
rect 338672 303340 338724 303346
rect 338672 303282 338724 303288
rect 338580 303068 338632 303074
rect 338580 303010 338632 303016
rect 338580 302388 338632 302394
rect 338580 302330 338632 302336
rect 338592 247586 338620 302330
rect 338868 300422 338896 310420
rect 339052 307873 339080 310420
rect 339038 307864 339094 307873
rect 339038 307799 339094 307808
rect 339236 306270 339264 310420
rect 339420 308582 339448 310420
rect 339408 308576 339460 308582
rect 339408 308518 339460 308524
rect 339604 308417 339632 310420
rect 339590 308408 339646 308417
rect 339590 308343 339646 308352
rect 339788 306354 339816 310420
rect 339972 308650 340000 310420
rect 339960 308644 340012 308650
rect 339960 308586 340012 308592
rect 340156 308553 340184 310420
rect 340142 308544 340198 308553
rect 340142 308479 340198 308488
rect 339604 306326 339816 306354
rect 339224 306264 339276 306270
rect 339224 306206 339276 306212
rect 338856 300416 338908 300422
rect 338856 300358 338908 300364
rect 339604 251122 339632 306326
rect 339684 306264 339736 306270
rect 339684 306206 339736 306212
rect 339696 300354 339724 306206
rect 339684 300348 339736 300354
rect 339684 300290 339736 300296
rect 340340 296714 340368 310420
rect 340524 306270 340552 310420
rect 340708 308961 340736 310420
rect 340694 308952 340750 308961
rect 340694 308887 340750 308896
rect 340892 308292 340920 310420
rect 341076 308854 341104 310420
rect 341064 308848 341116 308854
rect 341260 308825 341288 310420
rect 341064 308790 341116 308796
rect 341246 308816 341302 308825
rect 341246 308751 341302 308760
rect 340892 308264 341196 308292
rect 341064 306400 341116 306406
rect 341064 306342 341116 306348
rect 340512 306264 340564 306270
rect 340512 306206 340564 306212
rect 339972 296686 340368 296714
rect 339592 251116 339644 251122
rect 339592 251058 339644 251064
rect 339972 251054 340000 296686
rect 339960 251048 340012 251054
rect 339960 250990 340012 250996
rect 341076 250306 341104 306342
rect 341168 250442 341196 308264
rect 341444 308258 341472 310420
rect 341352 308230 341472 308258
rect 341248 308100 341300 308106
rect 341248 308042 341300 308048
rect 341156 250436 341208 250442
rect 341156 250378 341208 250384
rect 341064 250300 341116 250306
rect 341064 250242 341116 250248
rect 338580 247580 338632 247586
rect 338580 247522 338632 247528
rect 338488 243772 338540 243778
rect 338488 243714 338540 243720
rect 335728 243704 335780 243710
rect 335728 243646 335780 243652
rect 341260 243574 341288 308042
rect 341352 306406 341380 308230
rect 341432 308168 341484 308174
rect 341432 308110 341484 308116
rect 341340 306400 341392 306406
rect 341340 306342 341392 306348
rect 341444 248198 341472 308110
rect 341628 300490 341656 310420
rect 341812 308990 341840 310420
rect 341800 308984 341852 308990
rect 341800 308926 341852 308932
rect 341996 308106 342024 310420
rect 342180 308174 342208 310420
rect 342364 309126 342392 310420
rect 342352 309120 342404 309126
rect 342352 309062 342404 309068
rect 342352 308508 342404 308514
rect 342352 308450 342404 308456
rect 342168 308168 342220 308174
rect 342168 308110 342220 308116
rect 341984 308100 342036 308106
rect 341984 308042 342036 308048
rect 341616 300484 341668 300490
rect 341616 300426 341668 300432
rect 341432 248192 341484 248198
rect 341432 248134 341484 248140
rect 342364 247654 342392 308450
rect 342548 308394 342576 310420
rect 342732 308394 342760 310420
rect 342456 308366 342576 308394
rect 342640 308366 342760 308394
rect 342456 250782 342484 308366
rect 342536 308304 342588 308310
rect 342536 308246 342588 308252
rect 342444 250776 342496 250782
rect 342444 250718 342496 250724
rect 342548 250714 342576 308246
rect 342536 250708 342588 250714
rect 342536 250650 342588 250656
rect 342352 247648 342404 247654
rect 342352 247590 342404 247596
rect 342640 243642 342668 308366
rect 342916 297634 342944 310420
rect 343100 308310 343128 310420
rect 343284 308514 343312 310420
rect 343272 308508 343324 308514
rect 343272 308450 343324 308456
rect 343088 308304 343140 308310
rect 343088 308246 343140 308252
rect 343468 308242 343496 310420
rect 343456 308236 343508 308242
rect 343456 308178 343508 308184
rect 343652 307970 343680 310420
rect 343836 308394 343864 310420
rect 343744 308366 343864 308394
rect 343640 307964 343692 307970
rect 343640 307906 343692 307912
rect 342904 297628 342956 297634
rect 342904 297570 342956 297576
rect 343744 246906 343772 308366
rect 344020 306105 344048 310420
rect 344100 308644 344152 308650
rect 344100 308586 344152 308592
rect 344006 306096 344062 306105
rect 344006 306031 344062 306040
rect 343732 246900 343784 246906
rect 343732 246842 343784 246848
rect 344112 246838 344140 308586
rect 344204 308582 344232 310420
rect 344192 308576 344244 308582
rect 344192 308518 344244 308524
rect 344388 307834 344416 310420
rect 344376 307828 344428 307834
rect 344376 307770 344428 307776
rect 344572 306066 344600 310420
rect 344756 308514 344784 310420
rect 344940 308650 344968 310420
rect 344928 308644 344980 308650
rect 344928 308586 344980 308592
rect 344744 308508 344796 308514
rect 344744 308450 344796 308456
rect 345124 308394 345152 310420
rect 345308 308854 345336 310420
rect 345296 308848 345348 308854
rect 345296 308790 345348 308796
rect 345032 308366 345152 308394
rect 345204 308372 345256 308378
rect 344560 306060 344612 306066
rect 344560 306002 344612 306008
rect 345032 305998 345060 308366
rect 345204 308314 345256 308320
rect 345112 308304 345164 308310
rect 345112 308246 345164 308252
rect 345020 305992 345072 305998
rect 345020 305934 345072 305940
rect 345124 305930 345152 308246
rect 345112 305924 345164 305930
rect 345112 305866 345164 305872
rect 345216 305862 345244 308314
rect 345204 305856 345256 305862
rect 345204 305798 345256 305804
rect 344100 246832 344152 246838
rect 344100 246774 344152 246780
rect 345492 246770 345520 310420
rect 345676 308378 345704 310420
rect 345860 308922 345888 310420
rect 345848 308916 345900 308922
rect 345848 308858 345900 308864
rect 345664 308372 345716 308378
rect 345664 308314 345716 308320
rect 346044 296714 346072 310420
rect 346228 308310 346256 310420
rect 346412 308786 346440 310420
rect 346400 308780 346452 308786
rect 346400 308722 346452 308728
rect 346492 308644 346544 308650
rect 346492 308586 346544 308592
rect 346216 308304 346268 308310
rect 346216 308246 346268 308252
rect 345584 296686 346072 296714
rect 345480 246764 345532 246770
rect 345480 246706 345532 246712
rect 345584 244866 345612 296686
rect 346504 248266 346532 308586
rect 346492 248260 346544 248266
rect 346492 248202 346544 248208
rect 346596 248130 346624 310420
rect 346676 308304 346728 308310
rect 346676 308246 346728 308252
rect 346688 248198 346716 308246
rect 346780 254590 346808 310420
rect 346964 308650 346992 310420
rect 347148 308718 347176 310420
rect 347136 308712 347188 308718
rect 347136 308654 347188 308660
rect 346952 308644 347004 308650
rect 346952 308586 347004 308592
rect 346952 308372 347004 308378
rect 346952 308314 347004 308320
rect 346768 254584 346820 254590
rect 346768 254526 346820 254532
rect 346676 248192 346728 248198
rect 346676 248134 346728 248140
rect 346584 248124 346636 248130
rect 346584 248066 346636 248072
rect 346964 246294 346992 308314
rect 347332 305794 347360 310420
rect 347516 308310 347544 310420
rect 347700 308378 347728 310420
rect 347884 308394 347912 310420
rect 348068 308786 348096 310420
rect 348056 308780 348108 308786
rect 348056 308722 348108 308728
rect 348252 308394 348280 310420
rect 347688 308372 347740 308378
rect 347688 308314 347740 308320
rect 347792 308366 347912 308394
rect 348056 308372 348108 308378
rect 347504 308304 347556 308310
rect 347504 308246 347556 308252
rect 347320 305788 347372 305794
rect 347320 305730 347372 305736
rect 347792 305726 347820 308366
rect 348056 308314 348108 308320
rect 348160 308366 348280 308394
rect 348436 308378 348464 310420
rect 348424 308372 348476 308378
rect 348068 308122 348096 308314
rect 347884 308094 348096 308122
rect 347780 305720 347832 305726
rect 347780 305662 347832 305668
rect 347884 305658 347912 308094
rect 347964 306400 348016 306406
rect 347964 306342 348016 306348
rect 347872 305652 347924 305658
rect 347872 305594 347924 305600
rect 347976 248130 348004 306342
rect 347964 248124 348016 248130
rect 347964 248066 348016 248072
rect 348160 246702 348188 308366
rect 348424 308314 348476 308320
rect 348240 308304 348292 308310
rect 348240 308246 348292 308252
rect 348252 248334 348280 308246
rect 348620 306474 348648 310420
rect 348804 308310 348832 310420
rect 348792 308304 348844 308310
rect 348792 308246 348844 308252
rect 348608 306468 348660 306474
rect 348608 306410 348660 306416
rect 348988 303142 349016 310420
rect 349172 308378 349200 310420
rect 349252 308644 349304 308650
rect 349252 308586 349304 308592
rect 349160 308372 349212 308378
rect 349160 308314 349212 308320
rect 348976 303136 349028 303142
rect 348976 303078 349028 303084
rect 349264 303006 349292 308586
rect 349356 308394 349384 310420
rect 349540 308650 349568 310420
rect 349528 308644 349580 308650
rect 349528 308586 349580 308592
rect 349356 308366 349568 308394
rect 349344 308304 349396 308310
rect 349344 308246 349396 308252
rect 349252 303000 349304 303006
rect 349252 302942 349304 302948
rect 349356 250782 349384 308246
rect 349436 308236 349488 308242
rect 349436 308178 349488 308184
rect 349448 250850 349476 308178
rect 349436 250844 349488 250850
rect 349436 250786 349488 250792
rect 349344 250776 349396 250782
rect 349344 250718 349396 250724
rect 348240 248328 348292 248334
rect 348240 248270 348292 248276
rect 349540 247042 349568 308366
rect 349620 308372 349672 308378
rect 349620 308314 349672 308320
rect 349632 250714 349660 308314
rect 349724 308310 349752 310420
rect 349908 309058 349936 310420
rect 349896 309052 349948 309058
rect 349896 308994 349948 309000
rect 349712 308304 349764 308310
rect 349712 308246 349764 308252
rect 350092 302938 350120 310420
rect 350172 308916 350224 308922
rect 350172 308858 350224 308864
rect 350184 308650 350212 308858
rect 350172 308644 350224 308650
rect 350172 308586 350224 308592
rect 350276 308242 350304 310420
rect 350264 308236 350316 308242
rect 350264 308178 350316 308184
rect 350460 308174 350488 310420
rect 350644 308990 350672 310420
rect 350632 308984 350684 308990
rect 350632 308926 350684 308932
rect 350448 308168 350500 308174
rect 350448 308110 350500 308116
rect 350080 302932 350132 302938
rect 350080 302874 350132 302880
rect 350828 296714 350856 310420
rect 350644 296686 350856 296714
rect 349620 250708 349672 250714
rect 349620 250650 349672 250656
rect 349528 247036 349580 247042
rect 349528 246978 349580 246984
rect 350644 246702 350672 296686
rect 360856 258738 360884 446218
rect 360936 443760 360988 443766
rect 360936 443702 360988 443708
rect 360948 431934 360976 443702
rect 360936 431928 360988 431934
rect 360936 431870 360988 431876
rect 362236 325650 362264 446354
rect 363604 446344 363656 446350
rect 363604 446286 363656 446292
rect 362224 325644 362276 325650
rect 362224 325586 362276 325592
rect 363616 260166 363644 446286
rect 373264 446140 373316 446146
rect 373264 446082 373316 446088
rect 367744 443692 367796 443698
rect 367744 443634 367796 443640
rect 364984 443624 365036 443630
rect 364984 443566 365036 443572
rect 364996 273222 365024 443566
rect 367756 379506 367784 443634
rect 367744 379500 367796 379506
rect 367744 379442 367796 379448
rect 364984 273216 365036 273222
rect 364984 273158 365036 273164
rect 363604 260160 363656 260166
rect 363604 260102 363656 260108
rect 360844 258732 360896 258738
rect 360844 258674 360896 258680
rect 373276 254590 373304 446082
rect 454684 445868 454736 445874
rect 454684 445810 454736 445816
rect 442264 443352 442316 443358
rect 442264 443294 442316 443300
rect 436836 308848 436888 308854
rect 436836 308790 436888 308796
rect 436744 271380 436796 271386
rect 436744 271322 436796 271328
rect 373264 254584 373316 254590
rect 373264 254526 373316 254532
rect 348148 246696 348200 246702
rect 348148 246638 348200 246644
rect 350632 246696 350684 246702
rect 350632 246638 350684 246644
rect 346952 246288 347004 246294
rect 346952 246230 347004 246236
rect 345572 244860 345624 244866
rect 345572 244802 345624 244808
rect 342628 243636 342680 243642
rect 342628 243578 342680 243584
rect 341248 243568 341300 243574
rect 341248 243510 341300 243516
rect 299386 196072 299442 196081
rect 299386 196007 299442 196016
rect 299296 159112 299348 159118
rect 299296 159054 299348 159060
rect 299204 158364 299256 158370
rect 299204 158306 299256 158312
rect 299296 155372 299348 155378
rect 299296 155314 299348 155320
rect 299308 154834 299336 155314
rect 299296 154828 299348 154834
rect 299296 154770 299348 154776
rect 299400 9042 299428 196007
rect 316130 159896 316186 159905
rect 316130 159831 316186 159840
rect 336002 159896 336058 159905
rect 336002 159831 336058 159840
rect 338486 159896 338542 159905
rect 338486 159831 338542 159840
rect 348238 159896 348294 159905
rect 348238 159831 348294 159840
rect 351918 159896 351974 159905
rect 351918 159831 351974 159840
rect 363510 159896 363566 159905
rect 363510 159831 363566 159840
rect 370962 159896 371018 159905
rect 370962 159831 371018 159840
rect 299480 159656 299532 159662
rect 299480 159598 299532 159604
rect 299388 9036 299440 9042
rect 299388 8978 299440 8984
rect 298744 4072 298796 4078
rect 298744 4014 298796 4020
rect 299492 2774 299520 159598
rect 302240 159588 302292 159594
rect 302240 159530 302292 159536
rect 299572 151156 299624 151162
rect 299572 151098 299624 151104
rect 299584 7614 299612 151098
rect 300860 148368 300912 148374
rect 300860 148310 300912 148316
rect 300872 16574 300900 148310
rect 302252 16574 302280 159530
rect 316038 158672 316094 158681
rect 316038 158607 316094 158616
rect 316052 157146 316080 158607
rect 316040 157140 316092 157146
rect 316040 157082 316092 157088
rect 306380 156732 306432 156738
rect 306380 156674 306432 156680
rect 305000 153876 305052 153882
rect 305000 153818 305052 153824
rect 303620 146940 303672 146946
rect 303620 146882 303672 146888
rect 303632 16574 303660 146882
rect 305012 16574 305040 153818
rect 300872 16546 301544 16574
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 299572 7608 299624 7614
rect 299572 7550 299624 7556
rect 300768 7608 300820 7614
rect 300768 7550 300820 7556
rect 299492 2746 299704 2774
rect 299676 480 299704 2746
rect 300780 480 300808 7550
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 156674
rect 313280 156664 313332 156670
rect 313280 156606 313332 156612
rect 309138 155272 309194 155281
rect 309138 155207 309194 155216
rect 307760 134564 307812 134570
rect 307760 134506 307812 134512
rect 307772 3330 307800 134506
rect 307852 51740 307904 51746
rect 307852 51682 307904 51688
rect 307864 16574 307892 51682
rect 309152 16574 309180 155207
rect 310520 152720 310572 152726
rect 310520 152662 310572 152668
rect 310532 16574 310560 152662
rect 313292 16574 313320 156606
rect 314660 149796 314712 149802
rect 314660 149738 314712 149744
rect 307864 16546 307984 16574
rect 309152 16546 309824 16574
rect 310532 16546 311480 16574
rect 313292 16546 313872 16574
rect 307760 3324 307812 3330
rect 307760 3266 307812 3272
rect 307956 480 307984 16546
rect 309048 3324 309100 3330
rect 309048 3266 309100 3272
rect 309060 480 309088 3266
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311452 480 311480 16546
rect 312176 14476 312228 14482
rect 312176 14418 312228 14424
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 14418
rect 313844 480 313872 16546
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 149738
rect 316144 142154 316172 159831
rect 336016 159526 336044 159831
rect 336004 159520 336056 159526
rect 336004 159462 336056 159468
rect 338500 159458 338528 159831
rect 338488 159452 338540 159458
rect 338488 159394 338540 159400
rect 348252 159390 348280 159831
rect 350998 159760 351054 159769
rect 350998 159695 351054 159704
rect 348240 159384 348292 159390
rect 348240 159326 348292 159332
rect 351012 159322 351040 159695
rect 351000 159316 351052 159322
rect 351000 159258 351052 159264
rect 340972 158704 341024 158710
rect 316958 158672 317014 158681
rect 316958 158607 317014 158616
rect 318154 158672 318210 158681
rect 318154 158607 318210 158616
rect 319442 158672 319498 158681
rect 319442 158607 319498 158616
rect 320546 158672 320602 158681
rect 320546 158607 320602 158616
rect 321650 158672 321706 158681
rect 321650 158607 321706 158616
rect 323122 158672 323178 158681
rect 323122 158607 323178 158616
rect 326434 158672 326490 158681
rect 326434 158607 326490 158616
rect 328274 158672 328330 158681
rect 328274 158607 328330 158616
rect 329930 158672 329986 158681
rect 329930 158607 329986 158616
rect 330574 158672 330630 158681
rect 330574 158607 330630 158616
rect 333426 158672 333482 158681
rect 333426 158607 333482 158616
rect 334530 158672 334586 158681
rect 334530 158607 334586 158616
rect 335634 158672 335690 158681
rect 335634 158607 335690 158616
rect 338118 158672 338174 158681
rect 338118 158607 338174 158616
rect 340970 158672 340972 158681
rect 341024 158672 341026 158681
rect 340970 158607 341026 158616
rect 343546 158672 343602 158681
rect 343546 158607 343602 158616
rect 343914 158672 343970 158681
rect 343914 158607 343970 158616
rect 345938 158672 345994 158681
rect 345938 158607 345940 158616
rect 316972 156806 317000 158607
rect 318168 158098 318196 158607
rect 318156 158092 318208 158098
rect 318156 158034 318208 158040
rect 319456 157962 319484 158607
rect 319444 157956 319496 157962
rect 319444 157898 319496 157904
rect 320560 157894 320588 158607
rect 321664 158030 321692 158607
rect 321652 158024 321704 158030
rect 321652 157966 321704 157972
rect 320548 157888 320600 157894
rect 320548 157830 320600 157836
rect 321560 157412 321612 157418
rect 321560 157354 321612 157360
rect 316960 156800 317012 156806
rect 316960 156742 317012 156748
rect 321572 155378 321600 157354
rect 323136 156602 323164 158607
rect 326448 158166 326476 158607
rect 328288 158438 328316 158607
rect 328276 158432 328328 158438
rect 328276 158374 328328 158380
rect 329944 158302 329972 158607
rect 329932 158296 329984 158302
rect 329932 158238 329984 158244
rect 330588 158234 330616 158607
rect 333440 158370 333468 158607
rect 333610 158400 333666 158409
rect 333428 158364 333480 158370
rect 333610 158335 333666 158344
rect 333428 158306 333480 158312
rect 330576 158228 330628 158234
rect 330576 158170 330628 158176
rect 326436 158160 326488 158166
rect 326436 158102 326488 158108
rect 324226 157856 324282 157865
rect 324226 157791 324282 157800
rect 323124 156596 323176 156602
rect 323124 156538 323176 156544
rect 324240 155514 324268 157791
rect 329748 157480 329800 157486
rect 325330 157448 325386 157457
rect 329748 157422 329800 157428
rect 325330 157383 325386 157392
rect 324228 155508 324280 155514
rect 324228 155450 324280 155456
rect 321560 155372 321612 155378
rect 321560 155314 321612 155320
rect 325344 154154 325372 157383
rect 329760 154426 329788 157422
rect 333624 157214 333652 158335
rect 333612 157208 333664 157214
rect 333612 157150 333664 157156
rect 334544 157078 334572 158607
rect 334532 157072 334584 157078
rect 334532 157014 334584 157020
rect 335648 157010 335676 158607
rect 336830 158400 336886 158409
rect 336830 158335 336886 158344
rect 335636 157004 335688 157010
rect 335636 156946 335688 156952
rect 336844 156874 336872 158335
rect 338132 156942 338160 158607
rect 343560 158506 343588 158607
rect 343548 158500 343600 158506
rect 343548 158442 343600 158448
rect 338210 158264 338266 158273
rect 338210 158199 338266 158208
rect 338120 156936 338172 156942
rect 338120 156878 338172 156884
rect 336832 156868 336884 156874
rect 336832 156810 336884 156816
rect 338224 155922 338252 158199
rect 339498 157992 339554 158001
rect 339498 157927 339554 157936
rect 342350 157992 342406 158001
rect 342350 157927 342406 157936
rect 338212 155916 338264 155922
rect 338212 155858 338264 155864
rect 339512 155854 339540 157927
rect 341062 157856 341118 157865
rect 341062 157791 341118 157800
rect 339500 155848 339552 155854
rect 339500 155790 339552 155796
rect 341076 155582 341104 157791
rect 342364 155718 342392 157927
rect 343928 157350 343956 158607
rect 345992 158607 345994 158616
rect 348698 158672 348754 158681
rect 348698 158607 348754 158616
rect 345940 158578 345992 158584
rect 346674 157992 346730 158001
rect 346674 157927 346730 157936
rect 345110 157856 345166 157865
rect 345110 157791 345166 157800
rect 346398 157856 346454 157865
rect 346398 157791 346454 157800
rect 343916 157344 343968 157350
rect 343916 157286 343968 157292
rect 342352 155712 342404 155718
rect 342352 155654 342404 155660
rect 345124 155650 345152 157791
rect 345112 155644 345164 155650
rect 345112 155586 345164 155592
rect 341064 155576 341116 155582
rect 341064 155518 341116 155524
rect 346412 155446 346440 157791
rect 346688 155786 346716 157927
rect 348712 157282 348740 158607
rect 349802 157448 349858 157457
rect 349802 157383 349858 157392
rect 350998 157448 351054 157457
rect 350998 157383 351054 157392
rect 348700 157276 348752 157282
rect 348700 157218 348752 157224
rect 346676 155780 346728 155786
rect 346676 155722 346728 155728
rect 346400 155440 346452 155446
rect 346400 155382 346452 155388
rect 329748 154420 329800 154426
rect 329748 154362 329800 154368
rect 349816 154290 349844 157383
rect 349804 154284 349856 154290
rect 349804 154226 349856 154232
rect 351012 154222 351040 157383
rect 351000 154216 351052 154222
rect 351000 154158 351052 154164
rect 325332 154148 325384 154154
rect 325332 154090 325384 154096
rect 331220 152652 331272 152658
rect 331220 152594 331272 152600
rect 317420 145580 317472 145586
rect 317420 145522 317472 145528
rect 316052 142126 316172 142154
rect 316052 1154 316080 142126
rect 317432 16574 317460 145522
rect 328460 144220 328512 144226
rect 328460 144162 328512 144168
rect 318800 133204 318852 133210
rect 318800 133146 318852 133152
rect 318812 16574 318840 133146
rect 322940 89072 322992 89078
rect 322940 89014 322992 89020
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 316224 6860 316276 6866
rect 316224 6802 316276 6808
rect 316040 1148 316092 1154
rect 316040 1090 316092 1096
rect 316236 480 316264 6802
rect 317328 1148 317380 1154
rect 317328 1090 317380 1096
rect 317340 480 317368 1090
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 322112 6792 322164 6798
rect 322112 6734 322164 6740
rect 320914 3224 320970 3233
rect 320914 3159 320970 3168
rect 320928 480 320956 3159
rect 322124 480 322152 6734
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 354 322980 89014
rect 325700 89004 325752 89010
rect 325700 88946 325752 88952
rect 324320 22772 324372 22778
rect 324320 22714 324372 22720
rect 324332 3330 324360 22714
rect 325712 16574 325740 88946
rect 328472 16574 328500 144162
rect 329840 18624 329892 18630
rect 329840 18566 329892 18572
rect 329852 16574 329880 18566
rect 325712 16546 326384 16574
rect 328472 16546 328776 16574
rect 329852 16546 330432 16574
rect 324412 5024 324464 5030
rect 324412 4966 324464 4972
rect 324320 3324 324372 3330
rect 324320 3266 324372 3272
rect 324424 480 324452 4966
rect 325608 3324 325660 3330
rect 325608 3266 325660 3272
rect 325620 480 325648 3266
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328000 5092 328052 5098
rect 328000 5034 328052 5040
rect 328012 480 328040 5034
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 16546
rect 330404 480 330432 16546
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 152594
rect 333980 151088 334032 151094
rect 333980 151030 334032 151036
rect 332600 142860 332652 142866
rect 332600 142802 332652 142808
rect 332612 3210 332640 142802
rect 332692 131776 332744 131782
rect 332692 131718 332744 131724
rect 332704 3330 332732 131718
rect 333992 16574 334020 151030
rect 340880 149728 340932 149734
rect 340880 149670 340932 149676
rect 335360 141432 335412 141438
rect 335360 141374 335412 141380
rect 335372 16574 335400 141374
rect 339500 140072 339552 140078
rect 339500 140014 339552 140020
rect 333992 16546 334664 16574
rect 335372 16546 336320 16574
rect 332692 3324 332744 3330
rect 332692 3266 332744 3272
rect 333888 3324 333940 3330
rect 333888 3266 333940 3272
rect 332612 3182 332732 3210
rect 332704 480 332732 3182
rect 333900 480 333928 3266
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336292 480 336320 16546
rect 337474 8800 337530 8809
rect 337474 8735 337530 8744
rect 337488 480 337516 8735
rect 338672 4140 338724 4146
rect 338672 4082 338724 4088
rect 338684 480 338712 4082
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 354 339540 140014
rect 340892 3330 340920 149670
rect 345018 148336 345074 148345
rect 345018 148271 345074 148280
rect 342260 138712 342312 138718
rect 342260 138654 342312 138660
rect 340972 130416 341024 130422
rect 340972 130358 341024 130364
rect 340880 3324 340932 3330
rect 340880 3266 340932 3272
rect 340984 480 341012 130358
rect 342272 16574 342300 138654
rect 345032 16574 345060 148271
rect 350540 129056 350592 129062
rect 350540 128998 350592 129004
rect 350552 16574 350580 128998
rect 351932 16574 351960 159831
rect 353574 159760 353630 159769
rect 353574 159695 353630 159704
rect 356058 159760 356114 159769
rect 356058 159695 356114 159704
rect 360934 159760 360990 159769
rect 360934 159695 360990 159704
rect 353588 159254 353616 159695
rect 353576 159248 353628 159254
rect 353576 159190 353628 159196
rect 356072 159186 356100 159695
rect 356060 159180 356112 159186
rect 356060 159122 356112 159128
rect 360948 159050 360976 159695
rect 363524 159118 363552 159831
rect 363512 159112 363564 159118
rect 363512 159054 363564 159060
rect 360936 159044 360988 159050
rect 360936 158986 360988 158992
rect 370976 158982 371004 159831
rect 373998 159624 374054 159633
rect 373998 159559 374054 159568
rect 370964 158976 371016 158982
rect 370964 158918 371016 158924
rect 368204 158908 368256 158914
rect 368204 158850 368256 158856
rect 358452 158840 358504 158846
rect 358452 158782 358504 158788
rect 358464 158681 358492 158782
rect 368216 158681 368244 158850
rect 373356 158772 373408 158778
rect 373356 158714 373408 158720
rect 373368 158681 373396 158714
rect 355230 158672 355286 158681
rect 355230 158607 355286 158616
rect 356978 158672 357034 158681
rect 356978 158607 357034 158616
rect 358450 158672 358506 158681
rect 358450 158607 358506 158616
rect 365810 158672 365866 158681
rect 365810 158607 365866 158616
rect 368202 158672 368258 158681
rect 368202 158607 368258 158616
rect 373354 158672 373410 158681
rect 373354 158607 373410 158616
rect 353298 158264 353354 158273
rect 353298 158199 353354 158208
rect 352194 157448 352250 157457
rect 352194 157383 352250 157392
rect 352208 154358 352236 157383
rect 353312 154494 353340 158199
rect 355244 157486 355272 158607
rect 355232 157480 355284 157486
rect 354402 157448 354458 157457
rect 355232 157422 355284 157428
rect 356992 157418 357020 158607
rect 365824 158574 365852 158607
rect 365812 158568 365864 158574
rect 365812 158510 365864 158516
rect 354402 157383 354458 157392
rect 356980 157412 357032 157418
rect 354416 154562 354444 157383
rect 356980 157354 357032 157360
rect 354404 154556 354456 154562
rect 354404 154498 354456 154504
rect 353300 154488 353352 154494
rect 353300 154430 353352 154436
rect 352196 154352 352248 154358
rect 352196 154294 352248 154300
rect 357440 152584 357492 152590
rect 357440 152526 357492 152532
rect 342272 16546 342944 16574
rect 345032 16546 345336 16574
rect 350552 16546 351224 16574
rect 351932 16546 352880 16574
rect 342168 3324 342220 3330
rect 342168 3266 342220 3272
rect 342180 480 342208 3266
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344560 9240 344612 9246
rect 344560 9182 344612 9188
rect 344572 480 344600 9182
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 348056 9172 348108 9178
rect 348056 9114 348108 9120
rect 346952 3392 347004 3398
rect 346952 3334 347004 3340
rect 346964 480 346992 3334
rect 348068 480 348096 9114
rect 350448 6724 350500 6730
rect 350448 6666 350500 6672
rect 349252 4888 349304 4894
rect 349252 4830 349304 4836
rect 349264 480 349292 4830
rect 350460 480 350488 6666
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352852 480 352880 16546
rect 355232 9104 355284 9110
rect 355232 9046 355284 9052
rect 354036 6656 354088 6662
rect 354036 6598 354088 6604
rect 354048 480 354076 6598
rect 355244 480 355272 9046
rect 356334 4040 356390 4049
rect 356334 3975 356390 3984
rect 356348 480 356376 3975
rect 357452 3398 357480 152526
rect 364614 9616 364670 9625
rect 364614 9551 364670 9560
rect 361120 7608 361172 7614
rect 361120 7550 361172 7556
rect 362314 7576 362370 7585
rect 357532 6588 357584 6594
rect 357532 6530 357584 6536
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 357544 480 357572 6530
rect 359924 4820 359976 4826
rect 359924 4762 359976 4768
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 359936 480 359964 4762
rect 361132 480 361160 7550
rect 362314 7511 362370 7520
rect 362328 480 362356 7511
rect 363510 4992 363566 5001
rect 363510 4927 363566 4936
rect 363524 480 363552 4927
rect 364628 480 364656 9551
rect 370594 9480 370650 9489
rect 370594 9415 370650 9424
rect 365812 6520 365864 6526
rect 365812 6462 365864 6468
rect 365824 480 365852 6462
rect 368202 4856 368258 4865
rect 368202 4791 368258 4800
rect 367006 3904 367062 3913
rect 367006 3839 367062 3848
rect 367020 480 367048 3839
rect 368216 480 368244 4791
rect 369400 4072 369452 4078
rect 369400 4014 369452 4020
rect 369412 480 369440 4014
rect 370608 480 370636 9415
rect 372894 6896 372950 6905
rect 372894 6831 372950 6840
rect 371698 6080 371754 6089
rect 371698 6015 371754 6024
rect 371712 480 371740 6015
rect 372908 480 372936 6831
rect 374012 1170 374040 159559
rect 376758 159488 376814 159497
rect 376758 159423 376814 159432
rect 376024 158704 376076 158710
rect 376022 158672 376024 158681
rect 376076 158672 376078 158681
rect 376022 158607 376078 158616
rect 374092 152516 374144 152522
rect 374092 152458 374144 152464
rect 374104 3398 374132 152458
rect 376772 16574 376800 159423
rect 378138 159352 378194 159361
rect 378138 159287 378194 159296
rect 378152 16574 378180 159287
rect 378598 158672 378654 158681
rect 378598 158607 378600 158616
rect 378652 158607 378654 158616
rect 380990 158672 381046 158681
rect 380990 158607 381046 158616
rect 383566 158672 383622 158681
rect 383566 158607 383622 158616
rect 385958 158672 386014 158681
rect 385958 158607 386014 158616
rect 388534 158672 388590 158681
rect 388534 158607 388590 158616
rect 391478 158672 391534 158681
rect 391478 158607 391534 158616
rect 394238 158672 394294 158681
rect 394238 158607 394294 158616
rect 395894 158672 395950 158681
rect 395894 158607 395950 158616
rect 398470 158672 398526 158681
rect 398470 158607 398526 158616
rect 401046 158672 401102 158681
rect 401046 158607 401102 158616
rect 403990 158672 404046 158681
rect 403990 158607 404046 158616
rect 406474 158672 406530 158681
rect 406474 158607 406530 158616
rect 378600 158578 378652 158584
rect 381004 158574 381032 158607
rect 380992 158568 381044 158574
rect 380992 158510 381044 158516
rect 383580 158506 383608 158607
rect 383568 158500 383620 158506
rect 383568 158442 383620 158448
rect 385972 158438 386000 158607
rect 385960 158432 386012 158438
rect 385960 158374 386012 158380
rect 388548 158370 388576 158607
rect 388536 158364 388588 158370
rect 388536 158306 388588 158312
rect 391492 158302 391520 158607
rect 391480 158296 391532 158302
rect 391480 158238 391532 158244
rect 394252 158234 394280 158607
rect 394240 158228 394292 158234
rect 394240 158170 394292 158176
rect 395908 158166 395936 158607
rect 395896 158160 395948 158166
rect 395896 158102 395948 158108
rect 398484 158098 398512 158607
rect 398472 158092 398524 158098
rect 398472 158034 398524 158040
rect 401060 158030 401088 158607
rect 401048 158024 401100 158030
rect 401048 157966 401100 157972
rect 404004 157962 404032 158607
rect 403992 157956 404044 157962
rect 403992 157898 404044 157904
rect 406488 157894 406516 158607
rect 406476 157888 406528 157894
rect 406476 157830 406528 157836
rect 380898 152416 380954 152425
rect 380898 152351 380954 152360
rect 379518 82104 379574 82113
rect 379518 82039 379574 82048
rect 376772 16546 377720 16574
rect 378152 16546 378456 16574
rect 376024 10328 376076 10334
rect 376024 10270 376076 10276
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 10270
rect 377692 480 377720 16546
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 82039
rect 380912 16574 380940 152351
rect 380912 16546 381216 16574
rect 381188 480 381216 16546
rect 394238 9344 394294 9353
rect 394238 9279 394294 9288
rect 382370 6760 382426 6769
rect 382370 6695 382426 6704
rect 382384 480 382412 6695
rect 385958 6624 386014 6633
rect 385958 6559 386014 6568
rect 384764 4004 384816 4010
rect 384764 3946 384816 3952
rect 383566 3632 383622 3641
rect 383566 3567 383622 3576
rect 383580 480 383608 3567
rect 384776 480 384804 3946
rect 385972 480 386000 6559
rect 389454 6488 389510 6497
rect 389454 6423 389510 6432
rect 388258 3768 388314 3777
rect 388258 3703 388314 3712
rect 387154 3496 387210 3505
rect 387154 3431 387210 3440
rect 387168 480 387196 3431
rect 388272 480 388300 3703
rect 389468 480 389496 6423
rect 393042 6352 393098 6361
rect 393042 6287 393098 6296
rect 391848 3936 391900 3942
rect 391848 3878 391900 3884
rect 390650 3360 390706 3369
rect 390650 3295 390706 3304
rect 390664 480 390692 3295
rect 391860 480 391888 3878
rect 393056 480 393084 6287
rect 394252 480 394280 9279
rect 401322 9208 401378 9217
rect 401322 9143 401378 9152
rect 397736 9036 397788 9042
rect 397736 8978 397788 8984
rect 396538 6216 396594 6225
rect 396538 6151 396594 6160
rect 395344 3868 395396 3874
rect 395344 3810 395396 3816
rect 395356 480 395384 3810
rect 396552 480 396580 6151
rect 397748 480 397776 8978
rect 400128 6452 400180 6458
rect 400128 6394 400180 6400
rect 398932 3800 398984 3806
rect 398932 3742 398984 3748
rect 398944 480 398972 3742
rect 400140 480 400168 6394
rect 401336 480 401364 9143
rect 404818 9072 404874 9081
rect 404818 9007 404874 9016
rect 403624 6384 403676 6390
rect 403624 6326 403676 6332
rect 402520 3732 402572 3738
rect 402520 3674 402572 3680
rect 402532 480 402560 3674
rect 403636 480 403664 6326
rect 404832 480 404860 9007
rect 414296 8968 414348 8974
rect 411902 8936 411958 8945
rect 414296 8910 414348 8916
rect 411902 8871 411958 8880
rect 410800 6316 410852 6322
rect 410800 6258 410852 6264
rect 408408 6248 408460 6254
rect 408408 6190 408460 6196
rect 407212 6180 407264 6186
rect 407212 6122 407264 6128
rect 406016 3596 406068 3602
rect 406016 3538 406068 3544
rect 406028 480 406056 3538
rect 407224 480 407252 6122
rect 408420 480 408448 6190
rect 409604 3664 409656 3670
rect 409604 3606 409656 3612
rect 409616 480 409644 3606
rect 410812 480 410840 6258
rect 411916 480 411944 8871
rect 413100 3528 413152 3534
rect 413100 3470 413152 3476
rect 413112 480 413140 3470
rect 414308 480 414336 8910
rect 429660 4140 429712 4146
rect 429660 4082 429712 4088
rect 427268 4072 427320 4078
rect 427268 4014 427320 4020
rect 426164 4004 426216 4010
rect 426164 3946 426216 3952
rect 423772 3936 423824 3942
rect 423772 3878 423824 3884
rect 422576 3800 422628 3806
rect 422576 3742 422628 3748
rect 421380 3732 421432 3738
rect 421380 3674 421432 3680
rect 420184 3664 420236 3670
rect 420184 3606 420236 3612
rect 418988 3596 419040 3602
rect 418988 3538 419040 3544
rect 417884 3528 417936 3534
rect 417884 3470 417936 3476
rect 416688 3460 416740 3466
rect 416688 3402 416740 3408
rect 415492 3392 415544 3398
rect 415492 3334 415544 3340
rect 415504 480 415532 3334
rect 416700 480 416728 3402
rect 417896 480 417924 3470
rect 419000 480 419028 3538
rect 420196 480 420224 3606
rect 421392 480 421420 3674
rect 422588 480 422616 3742
rect 423784 480 423812 3878
rect 424968 3868 425020 3874
rect 424968 3810 425020 3816
rect 424980 480 425008 3810
rect 426176 480 426204 3946
rect 427280 480 427308 4014
rect 428464 3392 428516 3398
rect 428464 3334 428516 3340
rect 428476 480 428504 3334
rect 429672 480 429700 4082
rect 433246 3768 433302 3777
rect 433246 3703 433302 3712
rect 430856 3324 430908 3330
rect 430856 3266 430908 3272
rect 430868 480 430896 3266
rect 432052 3256 432104 3262
rect 432052 3198 432104 3204
rect 432064 480 432092 3198
rect 433260 480 433288 3703
rect 435546 3496 435602 3505
rect 435546 3431 435602 3440
rect 434442 3360 434498 3369
rect 434442 3295 434498 3304
rect 434456 480 434484 3295
rect 435560 480 435588 3431
rect 436756 480 436784 271322
rect 436848 158574 436876 308790
rect 440608 308780 440660 308786
rect 440608 308722 440660 308728
rect 439596 308712 439648 308718
rect 439596 308654 439648 308660
rect 438124 308644 438176 308650
rect 438124 308586 438176 308592
rect 438032 308576 438084 308582
rect 438032 308518 438084 308524
rect 436928 248260 436980 248266
rect 436928 248202 436980 248208
rect 436836 158568 436888 158574
rect 436836 158510 436888 158516
rect 436940 158370 436968 248202
rect 437480 248056 437532 248062
rect 437480 247998 437532 248004
rect 436928 158364 436980 158370
rect 436928 158306 436980 158312
rect 437492 4010 437520 247998
rect 437572 247988 437624 247994
rect 437572 247930 437624 247936
rect 437480 4004 437532 4010
rect 437480 3946 437532 3952
rect 437584 3602 437612 247930
rect 437756 245608 437808 245614
rect 437756 245550 437808 245556
rect 437664 245472 437716 245478
rect 437664 245414 437716 245420
rect 437676 3942 437704 245414
rect 437664 3936 437716 3942
rect 437664 3878 437716 3884
rect 437572 3596 437624 3602
rect 437572 3538 437624 3544
rect 437768 3398 437796 245550
rect 437848 245540 437900 245546
rect 437848 245482 437900 245488
rect 437860 4078 437888 245482
rect 437940 245268 437992 245274
rect 437940 245210 437992 245216
rect 437952 16574 437980 245210
rect 438044 158710 438072 308518
rect 438032 158704 438084 158710
rect 438032 158646 438084 158652
rect 438136 158506 438164 308586
rect 439504 308508 439556 308514
rect 439504 308450 439556 308456
rect 438860 308440 438912 308446
rect 438860 308382 438912 308388
rect 438216 250844 438268 250850
rect 438216 250786 438268 250792
rect 438124 158500 438176 158506
rect 438124 158442 438176 158448
rect 438228 157962 438256 250786
rect 438308 248192 438360 248198
rect 438308 248134 438360 248140
rect 438320 158302 438348 248134
rect 438308 158296 438360 158302
rect 438308 158238 438360 158244
rect 438216 157956 438268 157962
rect 438216 157898 438268 157904
rect 437952 16546 438072 16574
rect 437848 4072 437900 4078
rect 437848 4014 437900 4020
rect 438044 3738 438072 16546
rect 438032 3732 438084 3738
rect 438032 3674 438084 3680
rect 438872 3670 438900 308382
rect 438952 247852 439004 247858
rect 438952 247794 439004 247800
rect 438964 3806 438992 247794
rect 439044 247716 439096 247722
rect 439044 247658 439096 247664
rect 438952 3800 439004 3806
rect 438952 3742 439004 3748
rect 438860 3664 438912 3670
rect 437938 3632 437994 3641
rect 438860 3606 438912 3612
rect 437938 3567 437994 3576
rect 437756 3392 437808 3398
rect 437756 3334 437808 3340
rect 437952 480 437980 3567
rect 439056 3466 439084 247658
rect 439320 245404 439372 245410
rect 439320 245346 439372 245352
rect 439136 245200 439188 245206
rect 439136 245142 439188 245148
rect 439148 3874 439176 245142
rect 439228 245132 439280 245138
rect 439228 245074 439280 245080
rect 439136 3868 439188 3874
rect 439136 3810 439188 3816
rect 439240 3534 439268 245074
rect 439228 3528 439280 3534
rect 439134 3496 439190 3505
rect 439044 3460 439096 3466
rect 439228 3470 439280 3476
rect 439134 3431 439190 3440
rect 439044 3402 439096 3408
rect 439148 480 439176 3431
rect 439332 3330 439360 245346
rect 439412 245336 439464 245342
rect 439412 245278 439464 245284
rect 439424 16574 439452 245278
rect 439516 158642 439544 308450
rect 439504 158636 439556 158642
rect 439504 158578 439556 158584
rect 439608 158438 439636 308654
rect 440240 301572 440292 301578
rect 440240 301514 440292 301520
rect 439688 246696 439740 246702
rect 439688 246638 439740 246644
rect 439596 158432 439648 158438
rect 439596 158374 439648 158380
rect 439700 157894 439728 246638
rect 439688 157888 439740 157894
rect 439688 157830 439740 157836
rect 439424 16546 439544 16574
rect 439320 3324 439372 3330
rect 439320 3266 439372 3272
rect 439516 3262 439544 16546
rect 440252 3346 440280 301514
rect 440332 287768 440384 287774
rect 440332 287710 440384 287716
rect 440344 3534 440372 287710
rect 440424 247920 440476 247926
rect 440424 247862 440476 247868
rect 440436 3777 440464 247862
rect 440516 247784 440568 247790
rect 440516 247726 440568 247732
rect 440528 4146 440556 247726
rect 440620 158234 440648 308722
rect 441712 250776 441764 250782
rect 441712 250718 441764 250724
rect 441618 248160 441674 248169
rect 441618 248095 441674 248104
rect 440608 158228 440660 158234
rect 440608 158170 440660 158176
rect 441632 16574 441660 248095
rect 441724 158030 441752 250718
rect 441804 250708 441856 250714
rect 441804 250650 441856 250656
rect 441816 158098 441844 250650
rect 441896 248124 441948 248130
rect 441896 248066 441948 248072
rect 441908 158166 441936 248066
rect 441896 158160 441948 158166
rect 441896 158102 441948 158108
rect 441804 158092 441856 158098
rect 441804 158034 441856 158040
rect 441712 158024 441764 158030
rect 441712 157966 441764 157972
rect 442276 113150 442304 443294
rect 454696 438190 454724 445810
rect 580264 445052 580316 445058
rect 580264 444994 580316 445000
rect 494704 444780 494756 444786
rect 494704 444722 494756 444728
rect 454684 438184 454736 438190
rect 454684 438126 454736 438132
rect 478144 307148 478196 307154
rect 478144 307090 478196 307096
rect 458822 305960 458878 305969
rect 458822 305895 458878 305904
rect 445022 303240 445078 303249
rect 445022 303175 445078 303184
rect 442356 286476 442408 286482
rect 442356 286418 442408 286424
rect 442264 113144 442316 113150
rect 442264 113086 442316 113092
rect 441632 16546 442304 16574
rect 440516 4140 440568 4146
rect 440516 4082 440568 4088
rect 440422 3768 440478 3777
rect 440422 3703 440478 3712
rect 440332 3528 440384 3534
rect 440332 3470 440384 3476
rect 441528 3528 441580 3534
rect 441528 3470 441580 3476
rect 442276 3482 442304 16546
rect 442368 3602 442396 286418
rect 444380 280900 444432 280906
rect 444380 280842 444432 280848
rect 443000 253224 443052 253230
rect 443000 253166 443052 253172
rect 443012 16574 443040 253166
rect 443012 16546 443408 16574
rect 442356 3596 442408 3602
rect 442356 3538 442408 3544
rect 440252 3318 440372 3346
rect 439504 3256 439556 3262
rect 439504 3198 439556 3204
rect 440344 480 440372 3318
rect 441540 480 441568 3470
rect 442276 3454 442672 3482
rect 442644 480 442672 3454
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 444392 6914 444420 280842
rect 445036 16574 445064 303175
rect 449900 300280 449952 300286
rect 449900 300222 449952 300228
rect 448520 286408 448572 286414
rect 448520 286350 448572 286356
rect 446404 279540 446456 279546
rect 446404 279482 446456 279488
rect 445760 249280 445812 249286
rect 445760 249222 445812 249228
rect 445036 16546 445156 16574
rect 444392 6886 445064 6914
rect 445036 480 445064 6886
rect 445128 3466 445156 16546
rect 445116 3460 445168 3466
rect 445116 3402 445168 3408
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 249222
rect 446416 3398 446444 279482
rect 447416 3596 447468 3602
rect 447416 3538 447468 3544
rect 446404 3392 446456 3398
rect 446404 3334 446456 3340
rect 447428 480 447456 3538
rect 448532 3346 448560 286350
rect 448612 246628 448664 246634
rect 448612 246570 448664 246576
rect 448624 3534 448652 246570
rect 449912 16574 449940 300222
rect 453304 294840 453356 294846
rect 453304 294782 453356 294788
rect 452660 282328 452712 282334
rect 452660 282270 452712 282276
rect 452672 16574 452700 282270
rect 449912 16546 450952 16574
rect 452672 16546 453252 16574
rect 448612 3528 448664 3534
rect 448612 3470 448664 3476
rect 449808 3528 449860 3534
rect 449808 3470 449860 3476
rect 448532 3318 448652 3346
rect 448624 480 448652 3318
rect 449820 480 449848 3470
rect 450924 480 450952 16546
rect 453224 3482 453252 16546
rect 453316 3602 453344 294782
rect 454040 285116 454092 285122
rect 454040 285058 454092 285064
rect 453304 3596 453356 3602
rect 453304 3538 453356 3544
rect 453224 3454 453344 3482
rect 452108 3392 452160 3398
rect 452108 3334 452160 3340
rect 452120 480 452148 3334
rect 453316 480 453344 3454
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454052 354 454080 285058
rect 457444 278112 457496 278118
rect 457444 278054 457496 278060
rect 456892 250640 456944 250646
rect 456892 250582 456944 250588
rect 455696 3596 455748 3602
rect 455696 3538 455748 3544
rect 455708 480 455736 3538
rect 456904 480 456932 250582
rect 457456 2990 457484 278054
rect 458836 3466 458864 305895
rect 462964 298852 463016 298858
rect 462964 298794 463016 298800
rect 460940 282260 460992 282266
rect 460940 282202 460992 282208
rect 460204 276752 460256 276758
rect 460204 276694 460256 276700
rect 459560 250572 459612 250578
rect 459560 250514 459612 250520
rect 459572 16574 459600 250514
rect 459572 16546 459968 16574
rect 458088 3460 458140 3466
rect 458088 3402 458140 3408
rect 458824 3460 458876 3466
rect 458824 3402 458876 3408
rect 457444 2984 457496 2990
rect 457444 2926 457496 2932
rect 458100 480 458128 3402
rect 459192 2984 459244 2990
rect 459192 2926 459244 2932
rect 459204 480 459232 2926
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 460216 3874 460244 276694
rect 460952 16574 460980 282202
rect 460952 16546 461624 16574
rect 460204 3868 460256 3874
rect 460204 3810 460256 3816
rect 461596 480 461624 16546
rect 462780 3868 462832 3874
rect 462780 3810 462832 3816
rect 462792 480 462820 3810
rect 462976 3534 463004 298794
rect 476764 291916 476816 291922
rect 476764 291858 476816 291864
rect 471244 285048 471296 285054
rect 471244 284990 471296 284996
rect 464344 275392 464396 275398
rect 464344 275334 464396 275340
rect 463700 245064 463752 245070
rect 463700 245006 463752 245012
rect 463712 16574 463740 245006
rect 463712 16546 464016 16574
rect 462964 3528 463016 3534
rect 462964 3470 463016 3476
rect 463988 480 464016 16546
rect 464356 3058 464384 275334
rect 467104 273964 467156 273970
rect 467104 273906 467156 273912
rect 466460 260364 466512 260370
rect 466460 260306 466512 260312
rect 466472 16574 466500 260306
rect 466472 16546 467052 16574
rect 465172 3528 465224 3534
rect 465172 3470 465224 3476
rect 467024 3482 467052 16546
rect 467116 3602 467144 273906
rect 470600 258936 470652 258942
rect 470600 258878 470652 258884
rect 467840 252000 467892 252006
rect 467840 251942 467892 251948
rect 467852 16574 467880 251942
rect 467852 16546 468248 16574
rect 467104 3596 467156 3602
rect 467104 3538 467156 3544
rect 464344 3052 464396 3058
rect 464344 2994 464396 3000
rect 465184 480 465212 3470
rect 467024 3454 467512 3482
rect 466276 3052 466328 3058
rect 466276 2994 466328 3000
rect 466288 480 466316 2994
rect 467484 480 467512 3454
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 469864 3596 469916 3602
rect 469864 3538 469916 3544
rect 469876 480 469904 3538
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 470612 354 470640 258878
rect 471256 3126 471284 284990
rect 471980 283688 472032 283694
rect 471980 283630 472032 283636
rect 471992 16574 472020 283630
rect 473452 283620 473504 283626
rect 473452 283562 473504 283568
rect 473464 16574 473492 283562
rect 475384 271312 475436 271318
rect 475384 271254 475436 271260
rect 474740 268728 474792 268734
rect 474740 268670 474792 268676
rect 474752 16574 474780 268670
rect 471992 16546 472296 16574
rect 473464 16546 474136 16574
rect 474752 16546 475332 16574
rect 471244 3120 471296 3126
rect 471244 3062 471296 3068
rect 472268 480 472296 16546
rect 473452 3120 473504 3126
rect 473452 3062 473504 3068
rect 473464 480 473492 3062
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475304 3482 475332 16546
rect 475396 3602 475424 271254
rect 475384 3596 475436 3602
rect 475384 3538 475436 3544
rect 475304 3454 475792 3482
rect 475764 480 475792 3454
rect 476776 3194 476804 291858
rect 477500 268660 477552 268666
rect 477500 268602 477552 268608
rect 477512 6914 477540 268602
rect 478156 16574 478184 307090
rect 489920 307080 489972 307086
rect 489920 307022 489972 307028
rect 485044 304360 485096 304366
rect 485044 304302 485096 304308
rect 481640 270020 481692 270026
rect 481640 269962 481692 269968
rect 478156 16546 478276 16574
rect 477512 6886 478184 6914
rect 476948 3596 477000 3602
rect 476948 3538 477000 3544
rect 476764 3188 476816 3194
rect 476764 3130 476816 3136
rect 476960 480 476988 3538
rect 478156 480 478184 6886
rect 478248 3058 478276 16546
rect 481652 6914 481680 269962
rect 484400 268592 484452 268598
rect 484400 268534 484452 268540
rect 481732 249212 481784 249218
rect 481732 249154 481784 249160
rect 481744 16574 481772 249154
rect 484412 16574 484440 268534
rect 481744 16546 482416 16574
rect 484412 16546 484808 16574
rect 481652 6886 481772 6914
rect 479340 3188 479392 3194
rect 479340 3130 479392 3136
rect 478236 3052 478288 3058
rect 478236 2994 478288 3000
rect 479352 480 479380 3130
rect 480536 3052 480588 3058
rect 480536 2994 480588 3000
rect 480548 480 480576 2994
rect 481744 480 481772 6886
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484032 3460 484084 3466
rect 484032 3402 484084 3408
rect 484044 480 484072 3402
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 485056 3194 485084 304302
rect 485780 267164 485832 267170
rect 485780 267106 485832 267112
rect 485792 16574 485820 267106
rect 488540 258868 488592 258874
rect 488540 258810 488592 258816
rect 488552 16574 488580 258810
rect 485792 16546 486464 16574
rect 488552 16546 488856 16574
rect 485044 3188 485096 3194
rect 485044 3130 485096 3136
rect 486436 480 486464 16546
rect 487620 3188 487672 3194
rect 487620 3130 487672 3136
rect 487632 480 487660 3130
rect 488828 480 488856 16546
rect 489932 480 489960 307022
rect 494058 305824 494114 305833
rect 494058 305759 494114 305768
rect 492680 267096 492732 267102
rect 492680 267038 492732 267044
rect 491300 258800 491352 258806
rect 491300 258742 491352 258748
rect 490012 246560 490064 246566
rect 490012 246502 490064 246508
rect 490024 16574 490052 246502
rect 491312 16574 491340 258742
rect 492692 16574 492720 267038
rect 494072 16574 494100 305759
rect 494716 33114 494744 444722
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 579896 325644 579948 325650
rect 579896 325586 579948 325592
rect 579908 325281 579936 325586
rect 579894 325272 579950 325281
rect 579894 325207 579950 325216
rect 507860 304292 507912 304298
rect 507860 304234 507912 304240
rect 498290 303104 498346 303113
rect 498290 303039 498346 303048
rect 494796 267028 494848 267034
rect 494796 266970 494848 266976
rect 494704 33108 494756 33114
rect 494704 33050 494756 33056
rect 490024 16546 490696 16574
rect 491312 16546 492352 16574
rect 492692 16546 493088 16574
rect 494072 16546 494744 16574
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 492324 480 492352 16546
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 16546
rect 494716 480 494744 16546
rect 494808 2922 494836 266970
rect 496820 265736 496872 265742
rect 496820 265678 496872 265684
rect 495440 260296 495492 260302
rect 495440 260238 495492 260244
rect 494796 2916 494848 2922
rect 494796 2858 494848 2864
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 260238
rect 496832 16574 496860 265678
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498304 6914 498332 303039
rect 500224 301504 500276 301510
rect 500224 301446 500276 301452
rect 499580 279472 499632 279478
rect 499580 279414 499632 279420
rect 499592 16574 499620 279414
rect 499592 16546 500172 16574
rect 498212 6886 498332 6914
rect 498212 480 498240 6886
rect 500144 3482 500172 16546
rect 500236 3602 500264 301446
rect 502984 300212 503036 300218
rect 502984 300154 503036 300160
rect 502340 265668 502392 265674
rect 502340 265610 502392 265616
rect 502352 6914 502380 265610
rect 502996 16574 503024 300154
rect 504364 294772 504416 294778
rect 504364 294714 504416 294720
rect 503720 264376 503772 264382
rect 503720 264318 503772 264324
rect 502996 16546 503116 16574
rect 502352 6886 503024 6914
rect 500224 3596 500276 3602
rect 500224 3538 500276 3544
rect 501788 3596 501840 3602
rect 501788 3538 501840 3544
rect 500144 3454 500632 3482
rect 499396 2916 499448 2922
rect 499396 2858 499448 2864
rect 499408 480 499436 2858
rect 500604 480 500632 3454
rect 501800 480 501828 3538
rect 502996 480 503024 6886
rect 503088 3058 503116 16546
rect 503076 3052 503128 3058
rect 503076 2994 503128 3000
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 264318
rect 504376 3330 504404 294714
rect 506572 282192 506624 282198
rect 506572 282134 506624 282140
rect 506584 6914 506612 282134
rect 507872 16574 507900 304234
rect 514022 302968 514078 302977
rect 514022 302903 514078 302912
rect 512000 298784 512052 298790
rect 512000 298726 512052 298732
rect 509240 280832 509292 280838
rect 509240 280774 509292 280780
rect 509252 16574 509280 280774
rect 511264 264308 511316 264314
rect 511264 264250 511316 264256
rect 510620 263152 510672 263158
rect 510620 263094 510672 263100
rect 510632 16574 510660 263094
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 510632 16546 511212 16574
rect 506492 6886 506612 6914
rect 504364 3324 504416 3330
rect 504364 3266 504416 3272
rect 505376 3052 505428 3058
rect 505376 2994 505428 3000
rect 505388 480 505416 2994
rect 506492 480 506520 6886
rect 507676 3324 507728 3330
rect 507676 3266 507728 3272
rect 507688 480 507716 3266
rect 508884 480 508912 16546
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511184 3482 511212 16546
rect 511276 3602 511304 264250
rect 511264 3596 511316 3602
rect 511264 3538 511316 3544
rect 511184 3454 511304 3482
rect 511276 480 511304 3454
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 298726
rect 513564 3596 513616 3602
rect 513564 3538 513616 3544
rect 513576 480 513604 3538
rect 514036 3398 514064 302903
rect 561678 302832 561734 302841
rect 561678 302767 561734 302776
rect 554044 300144 554096 300150
rect 554044 300086 554096 300092
rect 516784 297424 516836 297430
rect 516784 297366 516836 297372
rect 516140 263084 516192 263090
rect 516140 263026 516192 263032
rect 514116 250504 514168 250510
rect 514116 250446 514168 250452
rect 514128 3466 514156 250446
rect 516152 16574 516180 263026
rect 516152 16546 516732 16574
rect 516704 3482 516732 16546
rect 516796 3874 516824 297366
rect 520924 296064 520976 296070
rect 520924 296006 520976 296012
rect 517520 278044 517572 278050
rect 517520 277986 517572 277992
rect 517532 16574 517560 277986
rect 520280 261724 520332 261730
rect 520280 261666 520332 261672
rect 517532 16546 517928 16574
rect 516784 3868 516836 3874
rect 516784 3810 516836 3816
rect 514116 3460 514168 3466
rect 514116 3402 514168 3408
rect 514760 3460 514812 3466
rect 516704 3454 517192 3482
rect 514760 3402 514812 3408
rect 514024 3392 514076 3398
rect 514024 3334 514076 3340
rect 514772 480 514800 3402
rect 515956 3392 516008 3398
rect 515956 3334 516008 3340
rect 515968 480 515996 3334
rect 517164 480 517192 3454
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 512430 -960 512542 326
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519544 3868 519596 3874
rect 519544 3810 519596 3816
rect 519556 480 519584 3810
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 261666
rect 520936 3126 520964 296006
rect 527824 294704 527876 294710
rect 527824 294646 527876 294652
rect 521660 276684 521712 276690
rect 521660 276626 521712 276632
rect 520924 3120 520976 3126
rect 520924 3062 520976 3068
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 276626
rect 524420 268524 524472 268530
rect 524420 268466 524472 268472
rect 523132 257372 523184 257378
rect 523132 257314 523184 257320
rect 523144 16574 523172 257314
rect 524432 16574 524460 268466
rect 527180 260228 527232 260234
rect 527180 260170 527232 260176
rect 525800 244996 525852 245002
rect 525800 244938 525852 244944
rect 525812 16574 525840 244938
rect 523144 16546 523816 16574
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 523040 3120 523092 3126
rect 523040 3062 523092 3068
rect 523052 480 523080 3062
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527192 6914 527220 260170
rect 527836 16574 527864 294646
rect 542360 294636 542412 294642
rect 542360 294578 542412 294584
rect 534724 293344 534776 293350
rect 534724 293286 534776 293292
rect 531320 261656 531372 261662
rect 531320 261598 531372 261604
rect 528560 251932 528612 251938
rect 528560 251874 528612 251880
rect 527836 16546 527956 16574
rect 527192 6886 527864 6914
rect 527836 480 527864 6886
rect 527928 3466 527956 16546
rect 527916 3460 527968 3466
rect 527916 3402 527968 3408
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 251874
rect 529938 248024 529994 248033
rect 529938 247959 529994 247968
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 247959
rect 531332 480 531360 261598
rect 531412 251864 531464 251870
rect 531412 251806 531464 251812
rect 531424 16574 531452 251806
rect 534078 247888 534134 247897
rect 534078 247823 534134 247832
rect 534092 16574 534120 247823
rect 531424 16546 532096 16574
rect 534092 16546 534488 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533712 3460 533764 3466
rect 533712 3402 533764 3408
rect 533724 480 533752 3402
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 534736 3194 534764 293286
rect 538864 291848 538916 291854
rect 538864 291790 538916 291796
rect 535460 261588 535512 261594
rect 535460 261530 535512 261536
rect 535472 16574 535500 261530
rect 538220 246492 538272 246498
rect 538220 246434 538272 246440
rect 535472 16546 536144 16574
rect 534724 3188 534776 3194
rect 534724 3130 534776 3136
rect 536116 480 536144 16546
rect 537208 3188 537260 3194
rect 537208 3130 537260 3136
rect 537220 480 537248 3130
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 246434
rect 538876 3534 538904 291790
rect 539692 275324 539744 275330
rect 539692 275266 539744 275272
rect 539704 6914 539732 275266
rect 540980 261520 541032 261526
rect 540980 261462 541032 261468
rect 540992 16574 541020 261462
rect 542372 16574 542400 294578
rect 553400 286340 553452 286346
rect 553400 286282 553452 286288
rect 546500 268456 546552 268462
rect 546500 268398 546552 268404
rect 545120 263016 545172 263022
rect 545120 262958 545172 262964
rect 543740 246424 543792 246430
rect 543740 246366 543792 246372
rect 543752 16574 543780 246366
rect 545132 16574 545160 262958
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 539612 6886 539732 6914
rect 538864 3528 538916 3534
rect 538864 3470 538916 3476
rect 539612 480 539640 6886
rect 540796 3528 540848 3534
rect 540796 3470 540848 3476
rect 540808 480 540836 3470
rect 542004 480 542032 16546
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 268398
rect 549260 268388 549312 268394
rect 549260 268330 549312 268336
rect 547880 262948 547932 262954
rect 547880 262890 547932 262896
rect 547892 3534 547920 262890
rect 547970 247752 548026 247761
rect 547970 247687 548026 247696
rect 547880 3528 547932 3534
rect 547880 3470 547932 3476
rect 547984 3346 548012 247687
rect 549272 16574 549300 268330
rect 552020 262880 552072 262886
rect 552020 262822 552072 262828
rect 550638 247616 550694 247625
rect 550638 247551 550694 247560
rect 550652 16574 550680 247551
rect 552032 16574 552060 262822
rect 553412 16574 553440 286282
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 548708 3528 548760 3534
rect 548708 3470 548760 3476
rect 547892 3318 548012 3346
rect 547892 480 547920 3318
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548720 354 548748 3470
rect 550284 480 550312 16546
rect 549046 354 549158 480
rect 548720 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 554056 3398 554084 300086
rect 560944 284980 560996 284986
rect 560944 284922 560996 284928
rect 560300 271244 560352 271250
rect 560300 271186 560352 271192
rect 556160 269952 556212 269958
rect 556160 269894 556212 269900
rect 554780 249144 554832 249150
rect 554780 249086 554832 249092
rect 554044 3392 554096 3398
rect 554044 3334 554096 3340
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 249086
rect 556172 3534 556200 269894
rect 556252 264240 556304 264246
rect 556252 264182 556304 264188
rect 556160 3528 556212 3534
rect 556160 3470 556212 3476
rect 556264 3346 556292 264182
rect 557540 249076 557592 249082
rect 557540 249018 557592 249024
rect 557552 16574 557580 249018
rect 560312 16574 560340 271186
rect 557552 16546 558592 16574
rect 560312 16546 560432 16574
rect 556988 3528 557040 3534
rect 556988 3470 557040 3476
rect 556172 3318 556292 3346
rect 556172 480 556200 3318
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557000 354 557028 3470
rect 558564 480 558592 16546
rect 559748 3392 559800 3398
rect 559748 3334 559800 3340
rect 559760 480 559788 3334
rect 557326 354 557438 480
rect 557000 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560404 354 560432 16546
rect 560956 3194 560984 284922
rect 561692 16574 561720 302767
rect 566464 295996 566516 296002
rect 566464 295938 566516 295944
rect 563704 290488 563756 290494
rect 563704 290430 563756 290436
rect 561692 16546 562088 16574
rect 560944 3188 560996 3194
rect 560944 3130 560996 3136
rect 562060 480 562088 16546
rect 563716 3534 563744 290430
rect 564532 246356 564584 246362
rect 564532 246298 564584 246304
rect 564544 6914 564572 246298
rect 565818 245168 565874 245177
rect 565818 245103 565874 245112
rect 565832 16574 565860 245103
rect 565832 16546 566412 16574
rect 564452 6886 564572 6914
rect 563704 3528 563756 3534
rect 563704 3470 563756 3476
rect 563244 3188 563296 3194
rect 563244 3130 563296 3136
rect 563256 480 563284 3130
rect 564452 480 564480 6886
rect 565636 3528 565688 3534
rect 565636 3470 565688 3476
rect 566384 3482 566412 16546
rect 566476 3874 566504 295938
rect 571340 293276 571392 293282
rect 571340 293218 571392 293224
rect 570604 289128 570656 289134
rect 570604 289070 570656 289076
rect 567844 271176 567896 271182
rect 567844 271118 567896 271124
rect 567200 269884 567252 269890
rect 567200 269826 567252 269832
rect 567212 16574 567240 269826
rect 567212 16546 567608 16574
rect 566464 3868 566516 3874
rect 566464 3810 566516 3816
rect 565648 480 565676 3470
rect 566384 3454 566872 3482
rect 566844 480 566872 3454
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567856 3194 567884 271118
rect 569132 3868 569184 3874
rect 569132 3810 569184 3816
rect 567844 3188 567896 3194
rect 567844 3130 567896 3136
rect 569144 480 569172 3810
rect 570616 3466 570644 289070
rect 570604 3460 570656 3466
rect 570604 3402 570656 3408
rect 570328 3188 570380 3194
rect 570328 3130 570380 3136
rect 570340 480 570368 3130
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 293218
rect 575480 287700 575532 287706
rect 575480 287642 575532 287648
rect 571984 269816 572036 269822
rect 571984 269758 572036 269764
rect 571996 3534 572024 269758
rect 574098 245032 574154 245041
rect 574098 244967 574154 244976
rect 574112 16574 574140 244967
rect 575492 16574 575520 287642
rect 579896 273216 579948 273222
rect 579896 273158 579948 273164
rect 579908 272241 579936 273158
rect 579894 272232 579950 272241
rect 579894 272167 579950 272176
rect 576860 244928 576912 244934
rect 576860 244870 576912 244876
rect 578238 244896 578294 244905
rect 576872 16574 576900 244870
rect 578238 244831 578294 244840
rect 578252 16574 578280 244831
rect 580276 152697 580304 444994
rect 581000 442264 581052 442270
rect 581000 442206 581052 442212
rect 580448 260160 580500 260166
rect 580448 260102 580500 260108
rect 580356 258732 580408 258738
rect 580356 258674 580408 258680
rect 580368 192545 580396 258674
rect 580460 232393 580488 260102
rect 580446 232384 580502 232393
rect 580446 232319 580502 232328
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 571984 3528 572036 3534
rect 571984 3470 572036 3476
rect 573916 3528 573968 3534
rect 573916 3470 573968 3476
rect 572720 3460 572772 3466
rect 572720 3402 572772 3408
rect 572732 480 572760 3402
rect 573928 480 573956 3470
rect 575124 480 575152 16546
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 581012 3534 581040 442206
rect 582380 438184 582432 438190
rect 582380 438126 582432 438132
rect 581092 254584 581144 254590
rect 581092 254526 581144 254532
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 581104 3346 581132 254526
rect 582392 16574 582420 438126
rect 582392 16546 583432 16574
rect 581828 3528 581880 3534
rect 581828 3470 581880 3476
rect 581012 3318 581132 3346
rect 581012 480 581040 3318
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 576278 -960 576390 326
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581840 354 581868 3470
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581840 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 3330 606056 3386 606112
rect 3330 579944 3386 580000
rect 3146 553832 3202 553888
rect 3330 527856 3386 527912
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 2870 501744 2926 501800
rect 3330 475632 3386 475688
rect 3330 462576 3386 462632
rect 2870 449520 2926 449576
rect 3514 658144 3570 658200
rect 3514 619112 3570 619168
rect 3606 566888 3662 566944
rect 217874 516840 217930 516896
rect 217782 515888 217838 515944
rect 217690 513712 217746 513768
rect 217598 489912 217654 489968
rect 217506 488280 217562 488336
rect 217322 488008 217378 488064
rect 219346 512760 219402 512816
rect 219162 510992 219218 511048
rect 219070 508136 219126 508192
rect 219254 509904 219310 509960
rect 242898 477264 242954 477320
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 3330 410488 3386 410544
rect 3330 397432 3386 397488
rect 3054 371320 3110 371376
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 3330 293120 3386 293176
rect 2962 267144 3018 267200
rect 3146 254088 3202 254144
rect 3238 241032 3294 241088
rect 3330 214920 3386 214976
rect 3146 188808 3202 188864
rect 3146 110608 3202 110664
rect 3606 358400 3662 358456
rect 3514 201864 3570 201920
rect 3514 162832 3570 162888
rect 3606 149776 3662 149832
rect 3514 136720 3570 136776
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 3422 45464 3478 45520
rect 3422 6432 3478 6488
rect 97906 305632 97962 305688
rect 97722 196832 97778 196888
rect 97814 195880 97870 195936
rect 97814 193704 97870 193760
rect 97722 192752 97778 192808
rect 97538 190984 97594 191040
rect 97446 188128 97502 188184
rect 97354 169904 97410 169960
rect 97630 189896 97686 189952
rect 97906 168408 97962 168464
rect 97906 168272 97962 168328
rect 230846 445712 230902 445768
rect 235906 476176 235962 476232
rect 237286 476332 237342 476368
rect 237286 476312 237288 476332
rect 237288 476312 237340 476332
rect 237340 476312 237342 476332
rect 237378 476176 237434 476232
rect 255226 476992 255282 477048
rect 264978 476992 265034 477048
rect 270498 476992 270554 477048
rect 304998 476992 305054 477048
rect 307758 476992 307814 477048
rect 244278 476604 244334 476640
rect 244278 476584 244280 476604
rect 244280 476584 244332 476604
rect 244332 476584 244334 476604
rect 247038 476584 247094 476640
rect 240230 476176 240286 476232
rect 241426 476176 241482 476232
rect 242806 476196 242862 476232
rect 244278 476312 244334 476368
rect 242806 476176 242808 476196
rect 242808 476176 242860 476196
rect 242860 476176 242862 476196
rect 245658 476176 245714 476232
rect 247222 476176 247278 476232
rect 249890 476448 249946 476504
rect 249798 476176 249854 476232
rect 255318 476856 255374 476912
rect 252558 476604 252614 476640
rect 252558 476584 252560 476604
rect 252560 476584 252612 476604
rect 252612 476584 252614 476604
rect 252466 476312 252522 476368
rect 251822 476176 251878 476232
rect 253202 476176 253258 476232
rect 254582 476176 254638 476232
rect 260838 476740 260894 476776
rect 260838 476720 260840 476740
rect 260840 476720 260892 476740
rect 260892 476720 260894 476740
rect 258078 476584 258134 476640
rect 258262 476584 258318 476640
rect 256606 476176 256662 476232
rect 257986 476176 258042 476232
rect 263598 476604 263654 476640
rect 263598 476584 263600 476604
rect 263600 476584 263652 476604
rect 263652 476584 263654 476604
rect 260746 476312 260802 476368
rect 261482 476176 261538 476232
rect 262126 476196 262182 476232
rect 262126 476176 262128 476196
rect 262128 476176 262180 476196
rect 262180 476176 262182 476196
rect 267922 476468 267978 476504
rect 267922 476448 267924 476468
rect 267924 476448 267976 476468
rect 267976 476448 267978 476468
rect 267646 476312 267702 476368
rect 263506 476176 263562 476232
rect 264886 476176 264942 476232
rect 266266 476176 266322 476232
rect 267554 476176 267610 476232
rect 277858 476856 277914 476912
rect 276018 476584 276074 476640
rect 273258 476448 273314 476504
rect 274454 476312 274510 476368
rect 269026 476176 269082 476232
rect 270406 476176 270462 476232
rect 271786 476176 271842 476232
rect 273166 476176 273222 476232
rect 274546 476176 274602 476232
rect 275926 476176 275982 476232
rect 277306 476176 277362 476232
rect 302238 476740 302294 476776
rect 302238 476720 302240 476740
rect 302240 476720 302292 476740
rect 302292 476720 302294 476740
rect 278686 476176 278742 476232
rect 280066 476176 280122 476232
rect 280250 476176 280306 476232
rect 283010 476176 283066 476232
rect 285770 476176 285826 476232
rect 287150 476176 287206 476232
rect 289910 476176 289966 476232
rect 292578 476176 292634 476232
rect 295430 476176 295486 476232
rect 298190 476176 298246 476232
rect 300858 476176 300914 476232
rect 297638 444352 297694 444408
rect 310518 476856 310574 476912
rect 313278 476448 313334 476504
rect 322938 476856 322994 476912
rect 314658 476468 314714 476504
rect 314658 476448 314660 476468
rect 314660 476448 314712 476468
rect 314712 476448 314714 476468
rect 317418 476332 317474 476368
rect 317418 476312 317420 476332
rect 317420 476312 317472 476332
rect 317472 476312 317474 476332
rect 320178 476312 320234 476368
rect 325790 476176 325846 476232
rect 580170 697176 580226 697232
rect 580262 683848 580318 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 579986 630808 580042 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 579894 537784 579950 537840
rect 580170 484608 580226 484664
rect 356518 445712 356574 445768
rect 158534 159840 158590 159896
rect 165986 159840 166042 159896
rect 173438 159840 173494 159896
rect 156050 159568 156106 159624
rect 206006 159568 206062 159624
rect 231858 159432 231914 159488
rect 213918 159296 213974 159352
rect 116490 158616 116546 158672
rect 117226 158616 117282 158672
rect 119710 158616 119766 158672
rect 120630 158652 120632 158672
rect 120632 158652 120684 158672
rect 120684 158652 120686 158672
rect 120630 158616 120686 158652
rect 121918 158616 121974 158672
rect 123206 158616 123262 158672
rect 126518 158616 126574 158672
rect 128174 158616 128230 158672
rect 128726 158616 128782 158672
rect 130566 158616 130622 158672
rect 131486 158616 131542 158672
rect 132406 158616 132462 158672
rect 133510 158616 133566 158672
rect 134890 158616 134946 158672
rect 158534 158616 158590 158672
rect 159914 158616 159970 158672
rect 160926 158616 160982 158672
rect 168286 158616 168342 158672
rect 118238 158344 118294 158400
rect 133694 158072 133750 158128
rect 124586 157528 124642 157584
rect 125414 157392 125470 157448
rect 135902 158480 135958 158536
rect 137006 158480 137062 158536
rect 138110 158480 138166 158536
rect 148874 158480 148930 158536
rect 136086 157800 136142 157856
rect 133694 155896 133750 155952
rect 141422 158208 141478 158264
rect 141790 158208 141846 158264
rect 144090 158208 144146 158264
rect 146022 158208 146078 158264
rect 146390 158208 146446 158264
rect 140686 157936 140742 157992
rect 140502 157800 140558 157856
rect 143078 157528 143134 157584
rect 145286 157800 145342 157856
rect 144366 157392 144422 157448
rect 144918 156576 144974 156632
rect 147678 157800 147734 157856
rect 148506 157392 148562 157448
rect 150990 158208 151046 158264
rect 149886 157392 149942 157448
rect 195886 158480 195942 158536
rect 178866 158344 178922 158400
rect 181810 158344 181866 158400
rect 184018 158344 184074 158400
rect 151358 157392 151414 157448
rect 152646 157392 152702 157448
rect 154118 157392 154174 157448
rect 154486 157392 154542 157448
rect 155774 157392 155830 157448
rect 157062 157392 157118 157448
rect 153198 155216 153254 155272
rect 175278 156712 175334 156768
rect 185950 158208 186006 158264
rect 178038 155352 178094 155408
rect 198462 157528 198518 157584
rect 201038 157528 201094 157584
rect 203430 157528 203486 157584
rect 202878 156848 202934 156904
rect 195978 152360 196034 152416
rect 220818 155488 220874 155544
rect 215298 138624 215354 138680
rect 222198 146920 222254 146976
rect 223578 127608 223634 127664
rect 238298 158072 238354 158128
rect 238482 157936 238538 157992
rect 240138 175888 240194 175944
rect 243542 308080 243598 308136
rect 256054 156712 256110 156768
rect 257802 308488 257858 308544
rect 257434 155216 257490 155272
rect 258262 3304 258318 3360
rect 261206 306448 261262 306504
rect 261482 306040 261538 306096
rect 261666 157256 261722 157312
rect 262678 156576 262734 156632
rect 264426 303456 264482 303512
rect 264426 155896 264482 155952
rect 265714 303320 265770 303376
rect 268290 155352 268346 155408
rect 268474 151000 268530 151056
rect 269854 158344 269910 158400
rect 270038 158208 270094 158264
rect 270590 308216 270646 308272
rect 270958 156848 271014 156904
rect 271602 158344 271658 158400
rect 271694 158208 271750 158264
rect 271418 157664 271474 157720
rect 273534 307944 273590 308000
rect 273350 307808 273406 307864
rect 274822 307944 274878 308000
rect 274638 307808 274694 307864
rect 273626 155488 273682 155544
rect 274454 158108 274456 158128
rect 274456 158108 274508 158128
rect 274508 158108 274510 158128
rect 274454 158072 274510 158108
rect 274362 157800 274418 157856
rect 274638 157548 274694 157584
rect 274638 157528 274640 157548
rect 274640 157528 274692 157548
rect 274692 157528 274694 157548
rect 275466 159432 275522 159488
rect 276018 158480 276074 158536
rect 275926 157528 275982 157584
rect 277030 158480 277086 158536
rect 277398 307808 277454 307864
rect 277950 158616 278006 158672
rect 278870 307808 278926 307864
rect 280158 307808 280214 307864
rect 280894 306040 280950 306096
rect 280894 157392 280950 157448
rect 283102 307808 283158 307864
rect 282182 125432 282238 125488
rect 283930 247016 283986 247072
rect 285034 247016 285090 247072
rect 286598 247016 286654 247072
rect 286966 158752 287022 158808
rect 288254 307808 288310 307864
rect 287794 247016 287850 247072
rect 288162 244296 288218 244352
rect 288346 158752 288402 158808
rect 289450 308896 289506 308952
rect 288990 159840 289046 159896
rect 289174 247016 289230 247072
rect 289726 158752 289782 158808
rect 290370 244704 290426 244760
rect 290646 158752 290702 158808
rect 290830 244432 290886 244488
rect 291106 244296 291162 244352
rect 291106 158752 291162 158808
rect 291750 244332 291752 244352
rect 291752 244332 291804 244352
rect 291804 244332 291806 244352
rect 291750 244296 291806 244332
rect 292486 308624 292542 308680
rect 292118 244296 292174 244352
rect 292486 158752 292542 158808
rect 292394 157392 292450 157448
rect 293774 307808 293830 307864
rect 293406 247016 293462 247072
rect 293406 244704 293462 244760
rect 293498 158752 293554 158808
rect 293774 245284 293776 245304
rect 293776 245284 293828 245304
rect 293828 245284 293830 245304
rect 293774 245248 293830 245284
rect 293774 245112 293830 245168
rect 293774 244296 293830 244352
rect 293774 167048 293830 167104
rect 293590 149096 293646 149152
rect 294326 159704 294382 159760
rect 295062 247052 295064 247072
rect 295064 247052 295116 247072
rect 295116 247052 295118 247072
rect 295062 247016 295118 247052
rect 294878 195200 294934 195256
rect 295246 244840 295302 244896
rect 295062 158752 295118 158808
rect 295798 245384 295854 245440
rect 295798 244840 295854 244896
rect 296350 307808 296406 307864
rect 296534 307808 296590 307864
rect 296626 244704 296682 244760
rect 296626 158752 296682 158808
rect 297270 308624 297326 308680
rect 298006 308080 298062 308136
rect 297822 307808 297878 307864
rect 296994 247968 297050 248024
rect 296902 247696 296958 247752
rect 297178 245112 297234 245168
rect 297362 244976 297418 245032
rect 297362 244432 297418 244488
rect 297270 196832 297326 196888
rect 297362 195880 297418 195936
rect 297454 193704 297510 193760
rect 297546 190984 297602 191040
rect 297362 189080 297418 189136
rect 297638 189896 297694 189952
rect 297638 189080 297694 189136
rect 297546 188128 297602 188184
rect 297638 169904 297694 169960
rect 297730 168000 297786 168056
rect 297914 168272 297970 168328
rect 298374 245520 298430 245576
rect 298282 159432 298338 159488
rect 298926 308080 298982 308136
rect 299110 307808 299166 307864
rect 298558 247288 298614 247344
rect 298466 159568 298522 159624
rect 299018 192752 299074 192808
rect 299110 188128 299166 188184
rect 299478 245384 299534 245440
rect 299754 245248 299810 245304
rect 299662 244840 299718 244896
rect 300122 248240 300178 248296
rect 300030 248104 300086 248160
rect 299938 247832 299994 247888
rect 299570 244568 299626 244624
rect 301226 245112 301282 245168
rect 301410 247424 301466 247480
rect 302514 247560 302570 247616
rect 303894 247288 303950 247344
rect 308310 297336 308366 297392
rect 308034 261432 308090 261488
rect 307942 248240 307998 248296
rect 307758 248104 307814 248160
rect 311254 303184 311310 303240
rect 306378 245248 306434 245304
rect 315394 305904 315450 305960
rect 316958 305768 317014 305824
rect 303802 244432 303858 244488
rect 301318 244296 301374 244352
rect 317970 303048 318026 303104
rect 320730 302912 320786 302968
rect 321650 247968 321706 248024
rect 324410 305632 324466 305688
rect 323030 247832 323086 247888
rect 325238 305632 325294 305688
rect 324410 247696 324466 247752
rect 325698 247560 325754 247616
rect 328090 302776 328146 302832
rect 327078 245112 327134 245168
rect 328458 244976 328514 245032
rect 330390 305496 330446 305552
rect 331310 308216 331366 308272
rect 330022 244840 330078 244896
rect 332230 306176 332286 306232
rect 333150 303456 333206 303512
rect 333978 303320 334034 303376
rect 339038 307808 339094 307864
rect 339590 308352 339646 308408
rect 340142 308488 340198 308544
rect 340694 308896 340750 308952
rect 341246 308760 341302 308816
rect 344006 306040 344062 306096
rect 299386 196016 299442 196072
rect 316130 159840 316186 159896
rect 336002 159840 336058 159896
rect 338486 159840 338542 159896
rect 348238 159840 348294 159896
rect 351918 159840 351974 159896
rect 363510 159840 363566 159896
rect 370962 159840 371018 159896
rect 316038 158616 316094 158672
rect 309138 155216 309194 155272
rect 350998 159704 351054 159760
rect 316958 158616 317014 158672
rect 318154 158616 318210 158672
rect 319442 158616 319498 158672
rect 320546 158616 320602 158672
rect 321650 158616 321706 158672
rect 323122 158616 323178 158672
rect 326434 158616 326490 158672
rect 328274 158616 328330 158672
rect 329930 158616 329986 158672
rect 330574 158616 330630 158672
rect 333426 158616 333482 158672
rect 334530 158616 334586 158672
rect 335634 158616 335690 158672
rect 338118 158616 338174 158672
rect 340970 158652 340972 158672
rect 340972 158652 341024 158672
rect 341024 158652 341026 158672
rect 340970 158616 341026 158652
rect 343546 158616 343602 158672
rect 343914 158616 343970 158672
rect 345938 158636 345994 158672
rect 345938 158616 345940 158636
rect 345940 158616 345992 158636
rect 345992 158616 345994 158636
rect 333610 158344 333666 158400
rect 324226 157800 324282 157856
rect 325330 157392 325386 157448
rect 336830 158344 336886 158400
rect 338210 158208 338266 158264
rect 339498 157936 339554 157992
rect 342350 157936 342406 157992
rect 341062 157800 341118 157856
rect 348698 158616 348754 158672
rect 346674 157936 346730 157992
rect 345110 157800 345166 157856
rect 346398 157800 346454 157856
rect 349802 157392 349858 157448
rect 350998 157392 351054 157448
rect 320914 3168 320970 3224
rect 337474 8744 337530 8800
rect 345018 148280 345074 148336
rect 353574 159704 353630 159760
rect 356058 159704 356114 159760
rect 360934 159704 360990 159760
rect 373998 159568 374054 159624
rect 355230 158616 355286 158672
rect 356978 158616 357034 158672
rect 358450 158616 358506 158672
rect 365810 158616 365866 158672
rect 368202 158616 368258 158672
rect 373354 158616 373410 158672
rect 353298 158208 353354 158264
rect 352194 157392 352250 157448
rect 354402 157392 354458 157448
rect 356334 3984 356390 4040
rect 364614 9560 364670 9616
rect 362314 7520 362370 7576
rect 363510 4936 363566 4992
rect 370594 9424 370650 9480
rect 368202 4800 368258 4856
rect 367006 3848 367062 3904
rect 372894 6840 372950 6896
rect 371698 6024 371754 6080
rect 376758 159432 376814 159488
rect 376022 158652 376024 158672
rect 376024 158652 376076 158672
rect 376076 158652 376078 158672
rect 376022 158616 376078 158652
rect 378138 159296 378194 159352
rect 378598 158636 378654 158672
rect 378598 158616 378600 158636
rect 378600 158616 378652 158636
rect 378652 158616 378654 158636
rect 380990 158616 381046 158672
rect 383566 158616 383622 158672
rect 385958 158616 386014 158672
rect 388534 158616 388590 158672
rect 391478 158616 391534 158672
rect 394238 158616 394294 158672
rect 395894 158616 395950 158672
rect 398470 158616 398526 158672
rect 401046 158616 401102 158672
rect 403990 158616 404046 158672
rect 406474 158616 406530 158672
rect 380898 152360 380954 152416
rect 379518 82048 379574 82104
rect 394238 9288 394294 9344
rect 382370 6704 382426 6760
rect 385958 6568 386014 6624
rect 383566 3576 383622 3632
rect 389454 6432 389510 6488
rect 388258 3712 388314 3768
rect 387154 3440 387210 3496
rect 393042 6296 393098 6352
rect 390650 3304 390706 3360
rect 401322 9152 401378 9208
rect 396538 6160 396594 6216
rect 404818 9016 404874 9072
rect 411902 8880 411958 8936
rect 433246 3712 433302 3768
rect 435546 3440 435602 3496
rect 434442 3304 434498 3360
rect 437938 3576 437994 3632
rect 439134 3440 439190 3496
rect 441618 248104 441674 248160
rect 458822 305904 458878 305960
rect 445022 303184 445078 303240
rect 440422 3712 440478 3768
rect 494058 305768 494114 305824
rect 580170 431568 580226 431624
rect 580170 378392 580226 378448
rect 579894 325216 579950 325272
rect 498290 303048 498346 303104
rect 514022 302912 514078 302968
rect 561678 302776 561734 302832
rect 529938 247968 529994 248024
rect 534078 247832 534134 247888
rect 547970 247696 548026 247752
rect 550638 247560 550694 247616
rect 565818 245112 565874 245168
rect 574098 244976 574154 245032
rect 579894 272176 579950 272232
rect 578238 244840 578294 244896
rect 580446 232328 580502 232384
rect 580354 192480 580410 192536
rect 580262 152632 580318 152688
rect 579802 112784 579858 112840
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
<< obsm2 >>
rect 220000 480000 356620 563308
rect 100000 160000 236620 243308
rect 300000 160000 436620 243308
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580257 683906 580323 683909
rect 583520 683906 584960 683996
rect 580257 683904 584960 683906
rect 580257 683848 580262 683904
rect 580318 683848 584960 683904
rect 580257 683846 584960 683848
rect 580257 683843 580323 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3325 606114 3391 606117
rect -960 606112 3391 606114
rect -960 606056 3330 606112
rect 3386 606056 3391 606112
rect -960 606054 3391 606056
rect -960 605964 480 606054
rect 3325 606051 3391 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3601 566946 3667 566949
rect -960 566944 3667 566946
rect -960 566888 3606 566944
rect 3662 566888 3667 566944
rect -960 566886 3667 566888
rect -960 566796 480 566886
rect 3601 566883 3667 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3141 553890 3207 553893
rect -960 553888 3207 553890
rect -960 553832 3146 553888
rect 3202 553832 3207 553888
rect -960 553830 3207 553832
rect -960 553740 480 553830
rect 3141 553827 3207 553830
rect -960 540684 480 540924
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 583520 551020 584960 551260
rect 579889 537842 579955 537845
rect 583520 537842 584960 537932
rect 579889 537840 584960 537842
rect 579889 537784 579894 537840
rect 579950 537784 584960 537840
rect 579889 537782 584960 537784
rect 579889 537779 579955 537782
rect 583520 537692 584960 537782
rect 583520 524364 584960 524604
rect 217869 516898 217935 516901
rect 219390 516898 220064 516924
rect 217869 516896 220064 516898
rect 217869 516840 217874 516896
rect 217930 516864 220064 516896
rect 217930 516840 219450 516864
rect 217869 516838 219450 516840
rect 217869 516835 217935 516838
rect 217777 515946 217843 515949
rect 219390 515946 220064 515972
rect 217777 515944 220064 515946
rect 217777 515888 217782 515944
rect 217838 515912 220064 515944
rect 217838 515888 219450 515912
rect 217777 515886 219450 515888
rect 217777 515883 217843 515886
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 217685 513770 217751 513773
rect 219390 513770 220064 513796
rect 217685 513768 220064 513770
rect 217685 513712 217690 513768
rect 217746 513736 220064 513768
rect 217746 513712 219450 513736
rect 217685 513710 219450 513712
rect 217685 513707 217751 513710
rect 219390 512821 220064 512844
rect 219341 512816 220064 512821
rect 219341 512760 219346 512816
rect 219402 512784 220064 512816
rect 219402 512760 219450 512784
rect 219341 512758 219450 512760
rect 219341 512755 219407 512758
rect 583520 511172 584960 511412
rect 219157 511050 219223 511053
rect 219390 511050 220064 511076
rect 219157 511048 220064 511050
rect 219157 510992 219162 511048
rect 219218 511016 220064 511048
rect 219218 510992 219450 511016
rect 219157 510990 219450 510992
rect 219157 510987 219223 510990
rect 219249 509962 219315 509965
rect 219390 509962 220064 509988
rect 219249 509960 220064 509962
rect 219249 509904 219254 509960
rect 219310 509928 220064 509960
rect 219310 509904 219450 509928
rect 219249 509902 219450 509904
rect 219249 509899 219315 509902
rect 219065 508194 219131 508197
rect 219390 508194 220064 508220
rect 219065 508192 220064 508194
rect 219065 508136 219070 508192
rect 219126 508160 220064 508192
rect 219126 508136 219450 508160
rect 219065 508134 219450 508136
rect 219065 508131 219131 508134
rect -960 501802 480 501892
rect 2865 501802 2931 501805
rect -960 501800 2931 501802
rect -960 501744 2870 501800
rect 2926 501744 2931 501800
rect -960 501742 2931 501744
rect -960 501652 480 501742
rect 2865 501739 2931 501742
rect 583520 497844 584960 498084
rect 217593 489970 217659 489973
rect 219390 489970 220064 489996
rect 217593 489968 220064 489970
rect 217593 489912 217598 489968
rect 217654 489936 220064 489968
rect 217654 489912 219450 489936
rect 217593 489910 219450 489912
rect 217593 489907 217659 489910
rect -960 488596 480 488836
rect 217501 488338 217567 488341
rect 219390 488338 220064 488364
rect 217501 488336 220064 488338
rect 217501 488280 217506 488336
rect 217562 488304 220064 488336
rect 217562 488280 219450 488304
rect 217501 488278 219450 488280
rect 217501 488275 217567 488278
rect 217317 488066 217383 488069
rect 219390 488066 220064 488092
rect 217317 488064 220064 488066
rect 217317 488008 217322 488064
rect 217378 488032 220064 488064
rect 217378 488008 219450 488032
rect 217317 488006 219450 488008
rect 217317 488003 217383 488006
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 242893 477322 242959 477325
rect 243118 477322 243124 477324
rect 242893 477320 243124 477322
rect 242893 477264 242898 477320
rect 242954 477264 243124 477320
rect 242893 477262 243124 477264
rect 242893 477259 242959 477262
rect 243118 477260 243124 477262
rect 243188 477260 243194 477324
rect 254526 476988 254532 477052
rect 254596 477050 254602 477052
rect 255221 477050 255287 477053
rect 254596 477048 255287 477050
rect 254596 476992 255226 477048
rect 255282 476992 255287 477048
rect 254596 476990 255287 476992
rect 254596 476988 254602 476990
rect 255221 476987 255287 476990
rect 264973 477050 265039 477053
rect 265934 477050 265940 477052
rect 264973 477048 265940 477050
rect 264973 476992 264978 477048
rect 265034 476992 265940 477048
rect 264973 476990 265940 476992
rect 264973 476987 265039 476990
rect 265934 476988 265940 476990
rect 266004 476988 266010 477052
rect 270493 477050 270559 477053
rect 270902 477050 270908 477052
rect 270493 477048 270908 477050
rect 270493 476992 270498 477048
rect 270554 476992 270908 477048
rect 270493 476990 270908 476992
rect 270493 476987 270559 476990
rect 270902 476988 270908 476990
rect 270972 476988 270978 477052
rect 304993 477050 305059 477053
rect 305862 477050 305868 477052
rect 304993 477048 305868 477050
rect 304993 476992 304998 477048
rect 305054 476992 305868 477048
rect 304993 476990 305868 476992
rect 304993 476987 305059 476990
rect 305862 476988 305868 476990
rect 305932 476988 305938 477052
rect 307753 477050 307819 477053
rect 308438 477050 308444 477052
rect 307753 477048 308444 477050
rect 307753 476992 307758 477048
rect 307814 476992 308444 477048
rect 307753 476990 308444 476992
rect 307753 476987 307819 476990
rect 308438 476988 308444 476990
rect 308508 476988 308514 477052
rect 255313 476914 255379 476917
rect 256182 476914 256188 476916
rect 255313 476912 256188 476914
rect 255313 476856 255318 476912
rect 255374 476856 256188 476912
rect 255313 476854 256188 476856
rect 255313 476851 255379 476854
rect 256182 476852 256188 476854
rect 256252 476852 256258 476916
rect 277853 476914 277919 476917
rect 278446 476914 278452 476916
rect 277853 476912 278452 476914
rect 277853 476856 277858 476912
rect 277914 476856 278452 476912
rect 277853 476854 278452 476856
rect 277853 476851 277919 476854
rect 278446 476852 278452 476854
rect 278516 476852 278522 476916
rect 310513 476914 310579 476917
rect 311014 476914 311020 476916
rect 310513 476912 311020 476914
rect 310513 476856 310518 476912
rect 310574 476856 311020 476912
rect 310513 476854 311020 476856
rect 310513 476851 310579 476854
rect 311014 476852 311020 476854
rect 311084 476852 311090 476916
rect 322933 476914 322999 476917
rect 323342 476914 323348 476916
rect 322933 476912 323348 476914
rect 322933 476856 322938 476912
rect 322994 476856 323348 476912
rect 322933 476854 323348 476856
rect 322933 476851 322999 476854
rect 323342 476852 323348 476854
rect 323412 476852 323418 476916
rect 260833 476778 260899 476781
rect 260966 476778 260972 476780
rect 260833 476776 260972 476778
rect 260833 476720 260838 476776
rect 260894 476720 260972 476776
rect 260833 476718 260972 476720
rect 260833 476715 260899 476718
rect 260966 476716 260972 476718
rect 261036 476716 261042 476780
rect 302233 476778 302299 476781
rect 303470 476778 303476 476780
rect 302233 476776 303476 476778
rect 302233 476720 302238 476776
rect 302294 476720 303476 476776
rect 302233 476718 303476 476720
rect 302233 476715 302299 476718
rect 303470 476716 303476 476718
rect 303540 476716 303546 476780
rect 244273 476644 244339 476645
rect 244222 476580 244228 476644
rect 244292 476642 244339 476644
rect 247033 476642 247099 476645
rect 248270 476642 248276 476644
rect 244292 476640 244384 476642
rect 244334 476584 244384 476640
rect 244292 476582 244384 476584
rect 247033 476640 248276 476642
rect 247033 476584 247038 476640
rect 247094 476584 248276 476640
rect 247033 476582 248276 476584
rect 244292 476580 244339 476582
rect 244273 476579 244339 476580
rect 247033 476579 247099 476582
rect 248270 476580 248276 476582
rect 248340 476580 248346 476644
rect 252553 476642 252619 476645
rect 253606 476642 253612 476644
rect 252553 476640 253612 476642
rect 252553 476584 252558 476640
rect 252614 476584 253612 476640
rect 252553 476582 253612 476584
rect 252553 476579 252619 476582
rect 253606 476580 253612 476582
rect 253676 476580 253682 476644
rect 257838 476580 257844 476644
rect 257908 476642 257914 476644
rect 258073 476642 258139 476645
rect 257908 476640 258139 476642
rect 257908 476584 258078 476640
rect 258134 476584 258139 476640
rect 257908 476582 258139 476584
rect 257908 476580 257914 476582
rect 258073 476579 258139 476582
rect 258257 476642 258323 476645
rect 263593 476644 263659 476645
rect 258390 476642 258396 476644
rect 258257 476640 258396 476642
rect 258257 476584 258262 476640
rect 258318 476584 258396 476640
rect 258257 476582 258396 476584
rect 258257 476579 258323 476582
rect 258390 476580 258396 476582
rect 258460 476580 258466 476644
rect 263542 476580 263548 476644
rect 263612 476642 263659 476644
rect 276013 476644 276079 476645
rect 276013 476642 276060 476644
rect 263612 476640 263704 476642
rect 263654 476584 263704 476640
rect 263612 476582 263704 476584
rect 275968 476640 276060 476642
rect 275968 476584 276018 476640
rect 275968 476582 276060 476584
rect 263612 476580 263659 476582
rect 263593 476579 263659 476580
rect 276013 476580 276060 476582
rect 276124 476580 276130 476644
rect 276013 476579 276079 476580
rect 249885 476506 249951 476509
rect 250662 476506 250668 476508
rect 249885 476504 250668 476506
rect 249885 476448 249890 476504
rect 249946 476448 250668 476504
rect 249885 476446 250668 476448
rect 249885 476443 249951 476446
rect 250662 476444 250668 476446
rect 250732 476444 250738 476508
rect 267917 476506 267983 476509
rect 268326 476506 268332 476508
rect 267917 476504 268332 476506
rect 267917 476448 267922 476504
rect 267978 476448 268332 476504
rect 267917 476446 268332 476448
rect 267917 476443 267983 476446
rect 268326 476444 268332 476446
rect 268396 476444 268402 476508
rect 273253 476506 273319 476509
rect 273478 476506 273484 476508
rect 273253 476504 273484 476506
rect 273253 476448 273258 476504
rect 273314 476448 273484 476504
rect 273253 476446 273484 476448
rect 273253 476443 273319 476446
rect 273478 476444 273484 476446
rect 273548 476444 273554 476508
rect 313273 476506 313339 476509
rect 313406 476506 313412 476508
rect 313273 476504 313412 476506
rect 313273 476448 313278 476504
rect 313334 476448 313412 476504
rect 313273 476446 313412 476448
rect 313273 476443 313339 476446
rect 313406 476444 313412 476446
rect 313476 476444 313482 476508
rect 314653 476506 314719 476509
rect 315798 476506 315804 476508
rect 314653 476504 315804 476506
rect 314653 476448 314658 476504
rect 314714 476448 315804 476504
rect 314653 476446 315804 476448
rect 314653 476443 314719 476446
rect 315798 476444 315804 476446
rect 315868 476444 315874 476508
rect 237281 476372 237347 476373
rect 237230 476308 237236 476372
rect 237300 476370 237347 476372
rect 244273 476370 244339 476373
rect 245326 476370 245332 476372
rect 237300 476368 237392 476370
rect 237342 476312 237392 476368
rect 237300 476310 237392 476312
rect 244273 476368 245332 476370
rect 244273 476312 244278 476368
rect 244334 476312 245332 476368
rect 244273 476310 245332 476312
rect 237300 476308 237347 476310
rect 237281 476307 237347 476308
rect 244273 476307 244339 476310
rect 245326 476308 245332 476310
rect 245396 476308 245402 476372
rect 251398 476308 251404 476372
rect 251468 476370 251474 476372
rect 252461 476370 252527 476373
rect 251468 476368 252527 476370
rect 251468 476312 252466 476368
rect 252522 476312 252527 476368
rect 251468 476310 252527 476312
rect 251468 476308 251474 476310
rect 252461 476307 252527 476310
rect 260598 476308 260604 476372
rect 260668 476370 260674 476372
rect 260741 476370 260807 476373
rect 260668 476368 260807 476370
rect 260668 476312 260746 476368
rect 260802 476312 260807 476368
rect 260668 476310 260807 476312
rect 260668 476308 260674 476310
rect 260741 476307 260807 476310
rect 266486 476308 266492 476372
rect 266556 476370 266562 476372
rect 267641 476370 267707 476373
rect 266556 476368 267707 476370
rect 266556 476312 267646 476368
rect 267702 476312 267707 476368
rect 266556 476310 267707 476312
rect 266556 476308 266562 476310
rect 267641 476307 267707 476310
rect 273294 476308 273300 476372
rect 273364 476370 273370 476372
rect 274449 476370 274515 476373
rect 273364 476368 274515 476370
rect 273364 476312 274454 476368
rect 274510 476312 274515 476368
rect 273364 476310 274515 476312
rect 273364 476308 273370 476310
rect 274449 476307 274515 476310
rect 317413 476370 317479 476373
rect 318374 476370 318380 476372
rect 317413 476368 318380 476370
rect 317413 476312 317418 476368
rect 317474 476312 318380 476368
rect 317413 476310 318380 476312
rect 317413 476307 317479 476310
rect 318374 476308 318380 476310
rect 318444 476308 318450 476372
rect 320173 476370 320239 476373
rect 320950 476370 320956 476372
rect 320173 476368 320956 476370
rect 320173 476312 320178 476368
rect 320234 476312 320956 476368
rect 320173 476310 320956 476312
rect 320173 476307 320239 476310
rect 320950 476308 320956 476310
rect 321020 476308 321026 476372
rect 235901 476236 235967 476237
rect 235901 476234 235948 476236
rect 235856 476232 235948 476234
rect 235856 476176 235906 476232
rect 235856 476174 235948 476176
rect 235901 476172 235948 476174
rect 236012 476172 236018 476236
rect 237373 476234 237439 476237
rect 238150 476234 238156 476236
rect 237373 476232 238156 476234
rect 237373 476176 237378 476232
rect 237434 476176 238156 476232
rect 237373 476174 238156 476176
rect 235901 476171 235967 476172
rect 237373 476171 237439 476174
rect 238150 476172 238156 476174
rect 238220 476172 238226 476236
rect 239622 476172 239628 476236
rect 239692 476234 239698 476236
rect 240225 476234 240291 476237
rect 239692 476232 240291 476234
rect 239692 476176 240230 476232
rect 240286 476176 240291 476232
rect 239692 476174 240291 476176
rect 239692 476172 239698 476174
rect 240225 476171 240291 476174
rect 240542 476172 240548 476236
rect 240612 476234 240618 476236
rect 241421 476234 241487 476237
rect 240612 476232 241487 476234
rect 240612 476176 241426 476232
rect 241482 476176 241487 476232
rect 240612 476174 241487 476176
rect 240612 476172 240618 476174
rect 241421 476171 241487 476174
rect 241830 476172 241836 476236
rect 241900 476234 241906 476236
rect 242801 476234 242867 476237
rect 241900 476232 242867 476234
rect 241900 476176 242806 476232
rect 242862 476176 242867 476232
rect 241900 476174 242867 476176
rect 241900 476172 241906 476174
rect 242801 476171 242867 476174
rect 245653 476234 245719 476237
rect 246430 476234 246436 476236
rect 245653 476232 246436 476234
rect 245653 476176 245658 476232
rect 245714 476176 246436 476232
rect 245653 476174 246436 476176
rect 245653 476171 245719 476174
rect 246430 476172 246436 476174
rect 246500 476172 246506 476236
rect 247217 476234 247283 476237
rect 247534 476234 247540 476236
rect 247217 476232 247540 476234
rect 247217 476176 247222 476232
rect 247278 476176 247540 476232
rect 247217 476174 247540 476176
rect 247217 476171 247283 476174
rect 247534 476172 247540 476174
rect 247604 476172 247610 476236
rect 248638 476172 248644 476236
rect 248708 476234 248714 476236
rect 249793 476234 249859 476237
rect 248708 476232 249859 476234
rect 248708 476176 249798 476232
rect 249854 476176 249859 476232
rect 248708 476174 249859 476176
rect 248708 476172 248714 476174
rect 249793 476171 249859 476174
rect 250110 476172 250116 476236
rect 250180 476234 250186 476236
rect 251817 476234 251883 476237
rect 250180 476232 251883 476234
rect 250180 476176 251822 476232
rect 251878 476176 251883 476232
rect 250180 476174 251883 476176
rect 250180 476172 250186 476174
rect 251817 476171 251883 476174
rect 252318 476172 252324 476236
rect 252388 476234 252394 476236
rect 253197 476234 253263 476237
rect 252388 476232 253263 476234
rect 252388 476176 253202 476232
rect 253258 476176 253263 476232
rect 252388 476174 253263 476176
rect 252388 476172 252394 476174
rect 253197 476171 253263 476174
rect 253422 476172 253428 476236
rect 253492 476234 253498 476236
rect 254577 476234 254643 476237
rect 253492 476232 254643 476234
rect 253492 476176 254582 476232
rect 254638 476176 254643 476232
rect 253492 476174 254643 476176
rect 253492 476172 253498 476174
rect 254577 476171 254643 476174
rect 255814 476172 255820 476236
rect 255884 476234 255890 476236
rect 256601 476234 256667 476237
rect 255884 476232 256667 476234
rect 255884 476176 256606 476232
rect 256662 476176 256667 476232
rect 255884 476174 256667 476176
rect 255884 476172 255890 476174
rect 256601 476171 256667 476174
rect 257102 476172 257108 476236
rect 257172 476234 257178 476236
rect 257981 476234 258047 476237
rect 257172 476232 258047 476234
rect 257172 476176 257986 476232
rect 258042 476176 258047 476232
rect 257172 476174 258047 476176
rect 257172 476172 257178 476174
rect 257981 476171 258047 476174
rect 259494 476172 259500 476236
rect 259564 476234 259570 476236
rect 261477 476234 261543 476237
rect 259564 476232 261543 476234
rect 259564 476176 261482 476232
rect 261538 476176 261543 476232
rect 259564 476174 261543 476176
rect 259564 476172 259570 476174
rect 261477 476171 261543 476174
rect 261702 476172 261708 476236
rect 261772 476234 261778 476236
rect 262121 476234 262187 476237
rect 261772 476232 262187 476234
rect 261772 476176 262126 476232
rect 262182 476176 262187 476232
rect 261772 476174 262187 476176
rect 261772 476172 261778 476174
rect 262121 476171 262187 476174
rect 262806 476172 262812 476236
rect 262876 476234 262882 476236
rect 263501 476234 263567 476237
rect 262876 476232 263567 476234
rect 262876 476176 263506 476232
rect 263562 476176 263567 476232
rect 262876 476174 263567 476176
rect 262876 476172 262882 476174
rect 263501 476171 263567 476174
rect 263910 476172 263916 476236
rect 263980 476234 263986 476236
rect 264881 476234 264947 476237
rect 263980 476232 264947 476234
rect 263980 476176 264886 476232
rect 264942 476176 264947 476232
rect 263980 476174 264947 476176
rect 263980 476172 263986 476174
rect 264881 476171 264947 476174
rect 265382 476172 265388 476236
rect 265452 476234 265458 476236
rect 266261 476234 266327 476237
rect 267549 476236 267615 476237
rect 267549 476234 267596 476236
rect 265452 476232 266327 476234
rect 265452 476176 266266 476232
rect 266322 476176 266327 476232
rect 265452 476174 266327 476176
rect 267504 476232 267596 476234
rect 267504 476176 267554 476232
rect 267504 476174 267596 476176
rect 265452 476172 265458 476174
rect 266261 476171 266327 476174
rect 267549 476172 267596 476174
rect 267660 476172 267666 476236
rect 268694 476172 268700 476236
rect 268764 476234 268770 476236
rect 269021 476234 269087 476237
rect 268764 476232 269087 476234
rect 268764 476176 269026 476232
rect 269082 476176 269087 476232
rect 268764 476174 269087 476176
rect 268764 476172 268770 476174
rect 267549 476171 267615 476172
rect 269021 476171 269087 476174
rect 269798 476172 269804 476236
rect 269868 476234 269874 476236
rect 270401 476234 270467 476237
rect 269868 476232 270467 476234
rect 269868 476176 270406 476232
rect 270462 476176 270467 476232
rect 269868 476174 270467 476176
rect 269868 476172 269874 476174
rect 270401 476171 270467 476174
rect 271270 476172 271276 476236
rect 271340 476234 271346 476236
rect 271781 476234 271847 476237
rect 271340 476232 271847 476234
rect 271340 476176 271786 476232
rect 271842 476176 271847 476232
rect 271340 476174 271847 476176
rect 271340 476172 271346 476174
rect 271781 476171 271847 476174
rect 272190 476172 272196 476236
rect 272260 476234 272266 476236
rect 273161 476234 273227 476237
rect 272260 476232 273227 476234
rect 272260 476176 273166 476232
rect 273222 476176 273227 476232
rect 272260 476174 273227 476176
rect 272260 476172 272266 476174
rect 273161 476171 273227 476174
rect 274398 476172 274404 476236
rect 274468 476234 274474 476236
rect 274541 476234 274607 476237
rect 275921 476236 275987 476237
rect 274468 476232 274607 476234
rect 274468 476176 274546 476232
rect 274602 476176 274607 476232
rect 274468 476174 274607 476176
rect 274468 476172 274474 476174
rect 274541 476171 274607 476174
rect 275870 476172 275876 476236
rect 275940 476234 275987 476236
rect 275940 476232 276032 476234
rect 275982 476176 276032 476232
rect 275940 476174 276032 476176
rect 275940 476172 275987 476174
rect 276974 476172 276980 476236
rect 277044 476234 277050 476236
rect 277301 476234 277367 476237
rect 277044 476232 277367 476234
rect 277044 476176 277306 476232
rect 277362 476176 277367 476232
rect 277044 476174 277367 476176
rect 277044 476172 277050 476174
rect 275921 476171 275987 476172
rect 277301 476171 277367 476174
rect 278078 476172 278084 476236
rect 278148 476234 278154 476236
rect 278681 476234 278747 476237
rect 278148 476232 278747 476234
rect 278148 476176 278686 476232
rect 278742 476176 278747 476232
rect 278148 476174 278747 476176
rect 278148 476172 278154 476174
rect 278681 476171 278747 476174
rect 279182 476172 279188 476236
rect 279252 476234 279258 476236
rect 280061 476234 280127 476237
rect 279252 476232 280127 476234
rect 279252 476176 280066 476232
rect 280122 476176 280127 476232
rect 279252 476174 280127 476176
rect 279252 476172 279258 476174
rect 280061 476171 280127 476174
rect 280245 476234 280311 476237
rect 280838 476234 280844 476236
rect 280245 476232 280844 476234
rect 280245 476176 280250 476232
rect 280306 476176 280844 476232
rect 280245 476174 280844 476176
rect 280245 476171 280311 476174
rect 280838 476172 280844 476174
rect 280908 476172 280914 476236
rect 283005 476234 283071 476237
rect 283414 476234 283420 476236
rect 283005 476232 283420 476234
rect 283005 476176 283010 476232
rect 283066 476176 283420 476232
rect 283005 476174 283420 476176
rect 283005 476171 283071 476174
rect 283414 476172 283420 476174
rect 283484 476172 283490 476236
rect 285765 476234 285831 476237
rect 285990 476234 285996 476236
rect 285765 476232 285996 476234
rect 285765 476176 285770 476232
rect 285826 476176 285996 476232
rect 285765 476174 285996 476176
rect 285765 476171 285831 476174
rect 285990 476172 285996 476174
rect 286060 476172 286066 476236
rect 287145 476234 287211 476237
rect 288198 476234 288204 476236
rect 287145 476232 288204 476234
rect 287145 476176 287150 476232
rect 287206 476176 288204 476232
rect 287145 476174 288204 476176
rect 287145 476171 287211 476174
rect 288198 476172 288204 476174
rect 288268 476172 288274 476236
rect 289905 476234 289971 476237
rect 290958 476234 290964 476236
rect 289905 476232 290964 476234
rect 289905 476176 289910 476232
rect 289966 476176 290964 476232
rect 289905 476174 290964 476176
rect 289905 476171 289971 476174
rect 290958 476172 290964 476174
rect 291028 476172 291034 476236
rect 292573 476234 292639 476237
rect 293350 476234 293356 476236
rect 292573 476232 293356 476234
rect 292573 476176 292578 476232
rect 292634 476176 293356 476232
rect 292573 476174 293356 476176
rect 292573 476171 292639 476174
rect 293350 476172 293356 476174
rect 293420 476172 293426 476236
rect 295425 476234 295491 476237
rect 295926 476234 295932 476236
rect 295425 476232 295932 476234
rect 295425 476176 295430 476232
rect 295486 476176 295932 476232
rect 295425 476174 295932 476176
rect 295425 476171 295491 476174
rect 295926 476172 295932 476174
rect 295996 476172 296002 476236
rect 298185 476234 298251 476237
rect 300853 476236 300919 476237
rect 298502 476234 298508 476236
rect 298185 476232 298508 476234
rect 298185 476176 298190 476232
rect 298246 476176 298508 476232
rect 298185 476174 298508 476176
rect 298185 476171 298251 476174
rect 298502 476172 298508 476174
rect 298572 476172 298578 476236
rect 300853 476234 300900 476236
rect 300808 476232 300900 476234
rect 300808 476176 300858 476232
rect 300808 476174 300900 476176
rect 300853 476172 300900 476174
rect 300964 476172 300970 476236
rect 325785 476234 325851 476237
rect 325918 476234 325924 476236
rect 325785 476232 325924 476234
rect 325785 476176 325790 476232
rect 325846 476176 325924 476232
rect 325785 476174 325924 476176
rect 300853 476171 300919 476172
rect 325785 476171 325851 476174
rect 325918 476172 325924 476174
rect 325988 476172 325994 476236
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 583520 471324 584960 471564
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 583520 457996 584960 458236
rect -960 449578 480 449668
rect 2865 449578 2931 449581
rect -960 449576 2931 449578
rect -960 449520 2870 449576
rect 2926 449520 2931 449576
rect -960 449518 2931 449520
rect -960 449428 480 449518
rect 2865 449515 2931 449518
rect 230841 445770 230907 445773
rect 356513 445770 356579 445773
rect 230841 445768 356579 445770
rect 230841 445712 230846 445768
rect 230902 445712 356518 445768
rect 356574 445712 356579 445768
rect 230841 445710 356579 445712
rect 230841 445707 230907 445710
rect 356513 445707 356579 445710
rect 583520 444668 584960 444908
rect 297633 444410 297699 444413
rect 439446 444410 439452 444412
rect 297633 444408 439452 444410
rect 297633 444352 297638 444408
rect 297694 444352 439452 444408
rect 297633 444350 439452 444352
rect 297633 444347 297699 444350
rect 439446 444348 439452 444350
rect 439516 444348 439522 444412
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 583520 418148 584960 418388
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 583520 404820 584960 405060
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3049 371378 3115 371381
rect -960 371376 3115 371378
rect -960 371320 3054 371376
rect 3110 371320 3115 371376
rect -960 371318 3115 371320
rect -960 371228 480 371318
rect 3049 371315 3115 371318
rect 583520 364972 584960 365212
rect -960 358458 480 358548
rect 3601 358458 3667 358461
rect -960 358456 3667 358458
rect -960 358400 3606 358456
rect 3662 358400 3667 358456
rect -960 358398 3667 358400
rect -960 358308 480 358398
rect 3601 358395 3667 358398
rect 583520 351780 584960 352020
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579889 325274 579955 325277
rect 583520 325274 584960 325364
rect 579889 325272 584960 325274
rect 579889 325216 579894 325272
rect 579950 325216 584960 325272
rect 579889 325214 584960 325216
rect 579889 325211 579955 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 583520 311932 584960 312172
rect 289445 308954 289511 308957
rect 340689 308954 340755 308957
rect 289445 308952 340755 308954
rect 289445 308896 289450 308952
rect 289506 308896 340694 308952
rect 340750 308896 340755 308952
rect 289445 308894 340755 308896
rect 289445 308891 289511 308894
rect 340689 308891 340755 308894
rect 286174 308756 286180 308820
rect 286244 308818 286250 308820
rect 341241 308818 341307 308821
rect 286244 308816 341307 308818
rect 286244 308760 341246 308816
rect 341302 308760 341307 308816
rect 286244 308758 341307 308760
rect 286244 308756 286250 308758
rect 341241 308755 341307 308758
rect 292481 308684 292547 308685
rect 292430 308682 292436 308684
rect 292390 308622 292436 308682
rect 292500 308680 292547 308684
rect 292542 308624 292547 308680
rect 292430 308620 292436 308622
rect 292500 308620 292547 308624
rect 292481 308619 292547 308620
rect 297265 308682 297331 308685
rect 297950 308682 297956 308684
rect 297265 308680 297956 308682
rect 297265 308624 297270 308680
rect 297326 308624 297956 308680
rect 297265 308622 297956 308624
rect 297265 308619 297331 308622
rect 297950 308620 297956 308622
rect 298020 308620 298026 308684
rect 257797 308546 257863 308549
rect 340137 308546 340203 308549
rect 257797 308544 340203 308546
rect 257797 308488 257802 308544
rect 257858 308488 340142 308544
rect 340198 308488 340203 308544
rect 257797 308486 340203 308488
rect 257797 308483 257863 308486
rect 340137 308483 340203 308486
rect 339585 308410 339651 308413
rect 248370 308408 339651 308410
rect 248370 308352 339590 308408
rect 339646 308352 339651 308408
rect 248370 308350 339651 308352
rect 243537 308138 243603 308141
rect 248370 308138 248430 308350
rect 339585 308347 339651 308350
rect 270585 308276 270651 308277
rect 270534 308274 270540 308276
rect 270494 308214 270540 308274
rect 270604 308272 270651 308276
rect 270646 308216 270651 308272
rect 270534 308212 270540 308214
rect 270604 308212 270651 308216
rect 284702 308212 284708 308276
rect 284772 308274 284778 308276
rect 331305 308274 331371 308277
rect 284772 308272 331371 308274
rect 284772 308216 331310 308272
rect 331366 308216 331371 308272
rect 284772 308214 331371 308216
rect 284772 308212 284778 308214
rect 270585 308211 270651 308212
rect 331305 308211 331371 308214
rect 243537 308136 248430 308138
rect 243537 308080 243542 308136
rect 243598 308080 248430 308136
rect 243537 308078 248430 308080
rect 243537 308075 243603 308078
rect 297766 308076 297772 308140
rect 297836 308138 297842 308140
rect 298001 308138 298067 308141
rect 297836 308136 298067 308138
rect 297836 308080 298006 308136
rect 298062 308080 298067 308136
rect 297836 308078 298067 308080
rect 297836 308076 297842 308078
rect 298001 308075 298067 308078
rect 298318 308076 298324 308140
rect 298388 308138 298394 308140
rect 298921 308138 298987 308141
rect 298388 308136 298987 308138
rect 298388 308080 298926 308136
rect 298982 308080 298987 308136
rect 298388 308078 298987 308080
rect 298388 308076 298394 308078
rect 298921 308075 298987 308078
rect 273294 307940 273300 308004
rect 273364 308002 273370 308004
rect 273529 308002 273595 308005
rect 273364 308000 273595 308002
rect 273364 307944 273534 308000
rect 273590 307944 273595 308000
rect 273364 307942 273595 307944
rect 273364 307940 273370 307942
rect 273529 307939 273595 307942
rect 274582 307940 274588 308004
rect 274652 308002 274658 308004
rect 274817 308002 274883 308005
rect 274652 308000 274883 308002
rect 274652 307944 274822 308000
rect 274878 307944 274883 308000
rect 274652 307942 274883 307944
rect 274652 307940 274658 307942
rect 274817 307939 274883 307942
rect 283414 307940 283420 308004
rect 283484 308002 283490 308004
rect 283484 307942 302250 308002
rect 283484 307940 283490 307942
rect 273345 307866 273411 307869
rect 273478 307866 273484 307868
rect 273345 307864 273484 307866
rect 273345 307808 273350 307864
rect 273406 307808 273484 307864
rect 273345 307806 273484 307808
rect 273345 307803 273411 307806
rect 273478 307804 273484 307806
rect 273548 307804 273554 307868
rect 274633 307866 274699 307869
rect 277393 307868 277459 307869
rect 278865 307868 278931 307869
rect 274766 307866 274772 307868
rect 274633 307864 274772 307866
rect 274633 307808 274638 307864
rect 274694 307808 274772 307864
rect 274633 307806 274772 307808
rect 274633 307803 274699 307806
rect 274766 307804 274772 307806
rect 274836 307804 274842 307868
rect 277342 307866 277348 307868
rect 277302 307806 277348 307866
rect 277412 307864 277459 307868
rect 278814 307866 278820 307868
rect 277454 307808 277459 307864
rect 277342 307804 277348 307806
rect 277412 307804 277459 307808
rect 278774 307806 278820 307866
rect 278884 307864 278931 307868
rect 278926 307808 278931 307864
rect 278814 307804 278820 307806
rect 278884 307804 278931 307808
rect 277393 307803 277459 307804
rect 278865 307803 278931 307804
rect 280153 307866 280219 307869
rect 283097 307868 283163 307869
rect 280286 307866 280292 307868
rect 280153 307864 280292 307866
rect 280153 307808 280158 307864
rect 280214 307808 280292 307864
rect 280153 307806 280292 307808
rect 280153 307803 280219 307806
rect 280286 307804 280292 307806
rect 280356 307804 280362 307868
rect 283046 307866 283052 307868
rect 283006 307806 283052 307866
rect 283116 307864 283163 307868
rect 283158 307808 283163 307864
rect 283046 307804 283052 307806
rect 283116 307804 283163 307808
rect 287830 307804 287836 307868
rect 287900 307866 287906 307868
rect 288249 307866 288315 307869
rect 293769 307868 293835 307869
rect 296345 307868 296411 307869
rect 296529 307868 296595 307869
rect 293718 307866 293724 307868
rect 287900 307864 288315 307866
rect 287900 307808 288254 307864
rect 288310 307808 288315 307864
rect 287900 307806 288315 307808
rect 293678 307806 293724 307866
rect 293788 307864 293835 307868
rect 296294 307866 296300 307868
rect 293830 307808 293835 307864
rect 287900 307804 287906 307806
rect 283097 307803 283163 307804
rect 288249 307803 288315 307806
rect 293718 307804 293724 307806
rect 293788 307804 293835 307808
rect 296254 307806 296300 307866
rect 296364 307864 296411 307868
rect 296406 307808 296411 307864
rect 296294 307804 296300 307806
rect 296364 307804 296411 307808
rect 296478 307804 296484 307868
rect 296548 307866 296595 307868
rect 296548 307864 296640 307866
rect 296590 307808 296640 307864
rect 296548 307806 296640 307808
rect 296548 307804 296595 307806
rect 297582 307804 297588 307868
rect 297652 307866 297658 307868
rect 297817 307866 297883 307869
rect 297652 307864 297883 307866
rect 297652 307808 297822 307864
rect 297878 307808 297883 307864
rect 297652 307806 297883 307808
rect 297652 307804 297658 307806
rect 293769 307803 293835 307804
rect 296345 307803 296411 307804
rect 296529 307803 296595 307804
rect 297817 307803 297883 307806
rect 298502 307804 298508 307868
rect 298572 307866 298578 307868
rect 299105 307866 299171 307869
rect 298572 307864 299171 307866
rect 298572 307808 299110 307864
rect 299166 307808 299171 307864
rect 298572 307806 299171 307808
rect 302190 307866 302250 307942
rect 339033 307866 339099 307869
rect 302190 307864 339099 307866
rect 302190 307808 339038 307864
rect 339094 307808 339099 307864
rect 302190 307806 339099 307808
rect 298572 307804 298578 307806
rect 299105 307803 299171 307806
rect 339033 307803 339099 307806
rect 261201 306506 261267 306509
rect 261201 306504 261402 306506
rect 261201 306448 261206 306504
rect 261262 306448 261402 306504
rect 261201 306446 261402 306448
rect 261201 306443 261267 306446
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 261342 306098 261402 306446
rect 278630 306172 278636 306236
rect 278700 306234 278706 306236
rect 332225 306234 332291 306237
rect 278700 306232 332291 306234
rect 278700 306176 332230 306232
rect 332286 306176 332291 306232
rect 278700 306174 332291 306176
rect 278700 306172 278706 306174
rect 332225 306171 332291 306174
rect 261477 306098 261543 306101
rect 261342 306096 261543 306098
rect 261342 306040 261482 306096
rect 261538 306040 261543 306096
rect 261342 306038 261543 306040
rect 261477 306035 261543 306038
rect 280889 306098 280955 306101
rect 344001 306098 344067 306101
rect 280889 306096 344067 306098
rect 280889 306040 280894 306096
rect 280950 306040 344006 306096
rect 344062 306040 344067 306096
rect 280889 306038 344067 306040
rect 280889 306035 280955 306038
rect 344001 306035 344067 306038
rect 315389 305962 315455 305965
rect 458817 305962 458883 305965
rect 315389 305960 458883 305962
rect 315389 305904 315394 305960
rect 315450 305904 458822 305960
rect 458878 305904 458883 305960
rect 315389 305902 458883 305904
rect 315389 305899 315455 305902
rect 458817 305899 458883 305902
rect 316953 305826 317019 305829
rect 494053 305826 494119 305829
rect 316953 305824 494119 305826
rect 316953 305768 316958 305824
rect 317014 305768 494058 305824
rect 494114 305768 494119 305824
rect 316953 305766 494119 305768
rect 316953 305763 317019 305766
rect 494053 305763 494119 305766
rect 97901 305690 97967 305693
rect 324405 305690 324471 305693
rect 325233 305690 325299 305693
rect 97901 305688 311910 305690
rect 97901 305632 97906 305688
rect 97962 305632 311910 305688
rect 97901 305630 311910 305632
rect 97901 305627 97967 305630
rect 311850 305554 311910 305630
rect 324405 305688 325299 305690
rect 324405 305632 324410 305688
rect 324466 305632 325238 305688
rect 325294 305632 325299 305688
rect 324405 305630 325299 305632
rect 324405 305627 324471 305630
rect 325233 305627 325299 305630
rect 330385 305554 330451 305557
rect 311850 305552 330451 305554
rect 311850 305496 330390 305552
rect 330446 305496 330451 305552
rect 311850 305494 330451 305496
rect 330385 305491 330451 305494
rect 264421 303514 264487 303517
rect 333145 303514 333211 303517
rect 264421 303512 333211 303514
rect 264421 303456 264426 303512
rect 264482 303456 333150 303512
rect 333206 303456 333211 303512
rect 264421 303454 333211 303456
rect 264421 303451 264487 303454
rect 333145 303451 333211 303454
rect 265709 303378 265775 303381
rect 333973 303378 334039 303381
rect 265709 303376 334039 303378
rect 265709 303320 265714 303376
rect 265770 303320 333978 303376
rect 334034 303320 334039 303376
rect 265709 303318 334039 303320
rect 265709 303315 265775 303318
rect 333973 303315 334039 303318
rect 311249 303242 311315 303245
rect 445017 303242 445083 303245
rect 311249 303240 445083 303242
rect 311249 303184 311254 303240
rect 311310 303184 445022 303240
rect 445078 303184 445083 303240
rect 311249 303182 445083 303184
rect 311249 303179 311315 303182
rect 445017 303179 445083 303182
rect 317965 303106 318031 303109
rect 498285 303106 498351 303109
rect 317965 303104 498351 303106
rect 317965 303048 317970 303104
rect 318026 303048 498290 303104
rect 498346 303048 498351 303104
rect 317965 303046 498351 303048
rect 317965 303043 318031 303046
rect 498285 303043 498351 303046
rect 320725 302970 320791 302973
rect 514017 302970 514083 302973
rect 320725 302968 514083 302970
rect 320725 302912 320730 302968
rect 320786 302912 514022 302968
rect 514078 302912 514083 302968
rect 320725 302910 514083 302912
rect 320725 302907 320791 302910
rect 514017 302907 514083 302910
rect 328085 302834 328151 302837
rect 561673 302834 561739 302837
rect 328085 302832 561739 302834
rect 328085 302776 328090 302832
rect 328146 302776 561678 302832
rect 561734 302776 561739 302832
rect 328085 302774 561739 302776
rect 328085 302771 328151 302774
rect 561673 302771 561739 302774
rect 583520 298604 584960 298844
rect 308305 297394 308371 297397
rect 437422 297394 437428 297396
rect 308305 297392 437428 297394
rect 308305 297336 308310 297392
rect 308366 297336 437428 297392
rect 308305 297334 437428 297336
rect 308305 297331 308371 297334
rect 437422 297332 437428 297334
rect 437492 297332 437498 297396
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579889 272234 579955 272237
rect 583520 272234 584960 272324
rect 579889 272232 584960 272234
rect 579889 272176 579894 272232
rect 579950 272176 584960 272232
rect 579889 272174 584960 272176
rect 579889 272171 579955 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2957 267202 3023 267205
rect -960 267200 3023 267202
rect -960 267144 2962 267200
rect 3018 267144 3023 267200
rect -960 267142 3023 267144
rect -960 267052 480 267142
rect 2957 267139 3023 267142
rect 308029 261490 308095 261493
rect 439078 261490 439084 261492
rect 308029 261488 439084 261490
rect 308029 261432 308034 261488
rect 308090 261432 439084 261488
rect 308029 261430 439084 261432
rect 308029 261427 308095 261430
rect 439078 261428 439084 261430
rect 439148 261428 439154 261492
rect 583520 258756 584960 258996
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 288198 248236 288204 248300
rect 288268 248298 288274 248300
rect 300117 248298 300183 248301
rect 288268 248296 300183 248298
rect 288268 248240 300122 248296
rect 300178 248240 300183 248296
rect 288268 248238 300183 248240
rect 288268 248236 288274 248238
rect 300117 248235 300183 248238
rect 307937 248298 308003 248301
rect 437606 248298 437612 248300
rect 307937 248296 437612 248298
rect 307937 248240 307942 248296
rect 307998 248240 437612 248296
rect 307937 248238 437612 248240
rect 307937 248235 308003 248238
rect 437606 248236 437612 248238
rect 437676 248236 437682 248300
rect 286910 248100 286916 248164
rect 286980 248162 286986 248164
rect 300025 248162 300091 248165
rect 286980 248160 300091 248162
rect 286980 248104 300030 248160
rect 300086 248104 300091 248160
rect 286980 248102 300091 248104
rect 286980 248100 286986 248102
rect 300025 248099 300091 248102
rect 307753 248162 307819 248165
rect 441613 248162 441679 248165
rect 307753 248160 441679 248162
rect 307753 248104 307758 248160
rect 307814 248104 441618 248160
rect 441674 248104 441679 248160
rect 307753 248102 441679 248104
rect 307753 248099 307819 248102
rect 441613 248099 441679 248102
rect 282310 247964 282316 248028
rect 282380 248026 282386 248028
rect 296989 248026 297055 248029
rect 282380 248024 297055 248026
rect 282380 247968 296994 248024
rect 297050 247968 297055 248024
rect 282380 247966 297055 247968
rect 282380 247964 282386 247966
rect 296989 247963 297055 247966
rect 321645 248026 321711 248029
rect 529933 248026 529999 248029
rect 321645 248024 529999 248026
rect 321645 247968 321650 248024
rect 321706 247968 529938 248024
rect 529994 247968 529999 248024
rect 321645 247966 529999 247968
rect 321645 247963 321711 247966
rect 529933 247963 529999 247966
rect 285070 247828 285076 247892
rect 285140 247890 285146 247892
rect 299933 247890 299999 247893
rect 285140 247888 299999 247890
rect 285140 247832 299938 247888
rect 299994 247832 299999 247888
rect 285140 247830 299999 247832
rect 285140 247828 285146 247830
rect 299933 247827 299999 247830
rect 323025 247890 323091 247893
rect 534073 247890 534139 247893
rect 323025 247888 534139 247890
rect 323025 247832 323030 247888
rect 323086 247832 534078 247888
rect 534134 247832 534139 247888
rect 323025 247830 534139 247832
rect 323025 247827 323091 247830
rect 534073 247827 534139 247830
rect 279918 247692 279924 247756
rect 279988 247754 279994 247756
rect 296897 247754 296963 247757
rect 279988 247752 296963 247754
rect 279988 247696 296902 247752
rect 296958 247696 296963 247752
rect 279988 247694 296963 247696
rect 279988 247692 279994 247694
rect 296897 247691 296963 247694
rect 324405 247754 324471 247757
rect 547965 247754 548031 247757
rect 324405 247752 548031 247754
rect 324405 247696 324410 247752
rect 324466 247696 547970 247752
rect 548026 247696 548031 247752
rect 324405 247694 548031 247696
rect 324405 247691 324471 247694
rect 547965 247691 548031 247694
rect 283966 247556 283972 247620
rect 284036 247618 284042 247620
rect 302509 247618 302575 247621
rect 284036 247616 302575 247618
rect 284036 247560 302514 247616
rect 302570 247560 302575 247616
rect 284036 247558 302575 247560
rect 284036 247556 284042 247558
rect 302509 247555 302575 247558
rect 325693 247618 325759 247621
rect 550633 247618 550699 247621
rect 325693 247616 550699 247618
rect 325693 247560 325698 247616
rect 325754 247560 550638 247616
rect 550694 247560 550699 247616
rect 325693 247558 550699 247560
rect 325693 247555 325759 247558
rect 550633 247555 550699 247558
rect 292246 247420 292252 247484
rect 292316 247482 292322 247484
rect 301405 247482 301471 247485
rect 292316 247480 301471 247482
rect 292316 247424 301410 247480
rect 301466 247424 301471 247480
rect 292316 247422 301471 247424
rect 292316 247420 292322 247422
rect 301405 247419 301471 247422
rect 298553 247346 298619 247349
rect 303889 247346 303955 247349
rect 298553 247344 303955 247346
rect 298553 247288 298558 247344
rect 298614 247288 303894 247344
rect 303950 247288 303955 247344
rect 298553 247286 303955 247288
rect 298553 247283 298619 247286
rect 303889 247283 303955 247286
rect 283925 247074 283991 247077
rect 284150 247074 284156 247076
rect 283925 247072 284156 247074
rect 283925 247016 283930 247072
rect 283986 247016 284156 247072
rect 283925 247014 284156 247016
rect 283925 247011 283991 247014
rect 284150 247012 284156 247014
rect 284220 247012 284226 247076
rect 284886 247012 284892 247076
rect 284956 247074 284962 247076
rect 285029 247074 285095 247077
rect 284956 247072 285095 247074
rect 284956 247016 285034 247072
rect 285090 247016 285095 247072
rect 284956 247014 285095 247016
rect 284956 247012 284962 247014
rect 285029 247011 285095 247014
rect 286358 247012 286364 247076
rect 286428 247074 286434 247076
rect 286593 247074 286659 247077
rect 286428 247072 286659 247074
rect 286428 247016 286598 247072
rect 286654 247016 286659 247072
rect 286428 247014 286659 247016
rect 286428 247012 286434 247014
rect 286593 247011 286659 247014
rect 287646 247012 287652 247076
rect 287716 247074 287722 247076
rect 287789 247074 287855 247077
rect 287716 247072 287855 247074
rect 287716 247016 287794 247072
rect 287850 247016 287855 247072
rect 287716 247014 287855 247016
rect 287716 247012 287722 247014
rect 287789 247011 287855 247014
rect 288750 247012 288756 247076
rect 288820 247074 288826 247076
rect 289169 247074 289235 247077
rect 288820 247072 289235 247074
rect 288820 247016 289174 247072
rect 289230 247016 289235 247072
rect 288820 247014 289235 247016
rect 288820 247012 288826 247014
rect 289169 247011 289235 247014
rect 293166 247012 293172 247076
rect 293236 247074 293242 247076
rect 293401 247074 293467 247077
rect 295057 247076 295123 247077
rect 295006 247074 295012 247076
rect 293236 247072 293467 247074
rect 293236 247016 293406 247072
rect 293462 247016 293467 247072
rect 293236 247014 293467 247016
rect 294966 247014 295012 247074
rect 295076 247072 295123 247076
rect 295118 247016 295123 247072
rect 293236 247012 293242 247014
rect 293401 247011 293467 247014
rect 295006 247012 295012 247014
rect 295076 247012 295123 247016
rect 295057 247011 295123 247012
rect 289302 245516 289308 245580
rect 289372 245578 289378 245580
rect 289372 245518 295994 245578
rect 289372 245516 289378 245518
rect 289118 245380 289124 245444
rect 289188 245442 289194 245444
rect 295793 245442 295859 245445
rect 289188 245440 295859 245442
rect 289188 245384 295798 245440
rect 295854 245384 295859 245440
rect 289188 245382 295859 245384
rect 289188 245380 289194 245382
rect 295793 245379 295859 245382
rect 293534 245244 293540 245308
rect 293604 245306 293610 245308
rect 293769 245306 293835 245309
rect 293604 245304 293835 245306
rect 293604 245248 293774 245304
rect 293830 245248 293835 245304
rect 293604 245246 293835 245248
rect 295934 245306 295994 245518
rect 298134 245516 298140 245580
rect 298204 245578 298210 245580
rect 298369 245578 298435 245581
rect 298204 245576 298435 245578
rect 298204 245520 298374 245576
rect 298430 245520 298435 245576
rect 298204 245518 298435 245520
rect 298204 245516 298210 245518
rect 298369 245515 298435 245518
rect 296110 245380 296116 245444
rect 296180 245442 296186 245444
rect 299473 245442 299539 245445
rect 296180 245440 299539 245442
rect 296180 245384 299478 245440
rect 299534 245384 299539 245440
rect 583520 245428 584960 245668
rect 296180 245382 299539 245384
rect 296180 245380 296186 245382
rect 299473 245379 299539 245382
rect 299749 245306 299815 245309
rect 295934 245304 299815 245306
rect 295934 245248 299754 245304
rect 299810 245248 299815 245304
rect 295934 245246 299815 245248
rect 293604 245244 293610 245246
rect 293769 245243 293835 245246
rect 299749 245243 299815 245246
rect 306373 245306 306439 245309
rect 437790 245306 437796 245308
rect 306373 245304 437796 245306
rect 306373 245248 306378 245304
rect 306434 245248 437796 245304
rect 306373 245246 437796 245248
rect 306373 245243 306439 245246
rect 437790 245244 437796 245246
rect 437860 245244 437866 245308
rect 286726 245108 286732 245172
rect 286796 245170 286802 245172
rect 293769 245170 293835 245173
rect 297173 245170 297239 245173
rect 286796 245168 293835 245170
rect 286796 245112 293774 245168
rect 293830 245112 293835 245168
rect 286796 245110 293835 245112
rect 286796 245108 286802 245110
rect 293769 245107 293835 245110
rect 294462 245168 297239 245170
rect 294462 245112 297178 245168
rect 297234 245112 297239 245168
rect 294462 245110 297239 245112
rect 282494 244972 282500 245036
rect 282564 245034 282570 245036
rect 294462 245034 294522 245110
rect 297173 245107 297239 245110
rect 299054 245108 299060 245172
rect 299124 245170 299130 245172
rect 301221 245170 301287 245173
rect 299124 245168 301287 245170
rect 299124 245112 301226 245168
rect 301282 245112 301287 245168
rect 299124 245110 301287 245112
rect 299124 245108 299130 245110
rect 301221 245107 301287 245110
rect 327073 245170 327139 245173
rect 565813 245170 565879 245173
rect 327073 245168 565879 245170
rect 327073 245112 327078 245168
rect 327134 245112 565818 245168
rect 565874 245112 565879 245168
rect 327073 245110 565879 245112
rect 327073 245107 327139 245110
rect 565813 245107 565879 245110
rect 297357 245034 297423 245037
rect 282564 244974 294522 245034
rect 294646 245032 297423 245034
rect 294646 244976 297362 245032
rect 297418 244976 297423 245032
rect 294646 244974 297423 244976
rect 282564 244972 282570 244974
rect 280470 244836 280476 244900
rect 280540 244898 280546 244900
rect 294646 244898 294706 244974
rect 297357 244971 297423 244974
rect 328453 245034 328519 245037
rect 574093 245034 574159 245037
rect 328453 245032 574159 245034
rect 328453 244976 328458 245032
rect 328514 244976 574098 245032
rect 574154 244976 574159 245032
rect 328453 244974 574159 244976
rect 328453 244971 328519 244974
rect 574093 244971 574159 244974
rect 295241 244900 295307 244901
rect 295190 244898 295196 244900
rect 280540 244838 294706 244898
rect 295150 244838 295196 244898
rect 295260 244896 295307 244900
rect 295302 244840 295307 244896
rect 280540 244836 280546 244838
rect 295190 244836 295196 244838
rect 295260 244836 295307 244840
rect 295241 244835 295307 244836
rect 295793 244898 295859 244901
rect 299657 244898 299723 244901
rect 295793 244896 299723 244898
rect 295793 244840 295798 244896
rect 295854 244840 299662 244896
rect 299718 244840 299723 244896
rect 295793 244838 299723 244840
rect 295793 244835 295859 244838
rect 299657 244835 299723 244838
rect 330017 244898 330083 244901
rect 578233 244898 578299 244901
rect 330017 244896 578299 244898
rect 330017 244840 330022 244896
rect 330078 244840 578238 244896
rect 578294 244840 578299 244896
rect 330017 244838 578299 244840
rect 330017 244835 330083 244838
rect 578233 244835 578299 244838
rect 282678 244700 282684 244764
rect 282748 244762 282754 244764
rect 290365 244762 290431 244765
rect 293401 244764 293467 244765
rect 293350 244762 293356 244764
rect 282748 244760 290431 244762
rect 282748 244704 290370 244760
rect 290426 244704 290431 244760
rect 282748 244702 290431 244704
rect 293310 244702 293356 244762
rect 293420 244760 293467 244764
rect 293462 244704 293467 244760
rect 282748 244700 282754 244702
rect 290365 244699 290431 244702
rect 293350 244700 293356 244702
rect 293420 244700 293467 244704
rect 295926 244700 295932 244764
rect 295996 244762 296002 244764
rect 296621 244762 296687 244765
rect 295996 244760 296687 244762
rect 295996 244704 296626 244760
rect 296682 244704 296687 244760
rect 295996 244702 296687 244704
rect 295996 244700 296002 244702
rect 293401 244699 293467 244700
rect 296621 244699 296687 244702
rect 289486 244564 289492 244628
rect 289556 244626 289562 244628
rect 299565 244626 299631 244629
rect 289556 244624 299631 244626
rect 289556 244568 299570 244624
rect 299626 244568 299631 244624
rect 289556 244566 299631 244568
rect 289556 244564 289562 244566
rect 299565 244563 299631 244566
rect 290825 244492 290891 244493
rect 290774 244490 290780 244492
rect 290734 244430 290780 244490
rect 290844 244488 290891 244492
rect 290886 244432 290891 244488
rect 290774 244428 290780 244430
rect 290844 244428 290891 244432
rect 290825 244427 290891 244428
rect 297357 244490 297423 244493
rect 303797 244490 303863 244493
rect 297357 244488 303863 244490
rect 297357 244432 297362 244488
rect 297418 244432 303802 244488
rect 303858 244432 303863 244488
rect 297357 244430 303863 244432
rect 297357 244427 297423 244430
rect 303797 244427 303863 244430
rect 288014 244292 288020 244356
rect 288084 244354 288090 244356
rect 288157 244354 288223 244357
rect 288084 244352 288223 244354
rect 288084 244296 288162 244352
rect 288218 244296 288223 244352
rect 288084 244294 288223 244296
rect 288084 244292 288090 244294
rect 288157 244291 288223 244294
rect 290590 244292 290596 244356
rect 290660 244354 290666 244356
rect 291101 244354 291167 244357
rect 291745 244356 291811 244357
rect 291694 244354 291700 244356
rect 290660 244352 291167 244354
rect 290660 244296 291106 244352
rect 291162 244296 291167 244352
rect 290660 244294 291167 244296
rect 291654 244294 291700 244354
rect 291764 244352 291811 244356
rect 291806 244296 291811 244352
rect 290660 244292 290666 244294
rect 291101 244291 291167 244294
rect 291694 244292 291700 244294
rect 291764 244292 291811 244296
rect 291878 244292 291884 244356
rect 291948 244354 291954 244356
rect 292113 244354 292179 244357
rect 291948 244352 292179 244354
rect 291948 244296 292118 244352
rect 292174 244296 292179 244352
rect 291948 244294 292179 244296
rect 291948 244292 291954 244294
rect 291745 244291 291811 244292
rect 292113 244291 292179 244294
rect 293769 244354 293835 244357
rect 301313 244354 301379 244357
rect 293769 244352 301379 244354
rect 293769 244296 293774 244352
rect 293830 244296 301318 244352
rect 301374 244296 301379 244352
rect 293769 244294 301379 244296
rect 293769 244291 293835 244294
rect 301313 244291 301379 244294
rect -960 241090 480 241180
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect -960 227884 480 228124
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect -960 201922 480 202012
rect 3509 201922 3575 201925
rect -960 201920 3575 201922
rect -960 201864 3514 201920
rect 3570 201864 3575 201920
rect -960 201862 3575 201864
rect -960 201772 480 201862
rect 3509 201859 3575 201862
rect 580441 232386 580507 232389
rect 583520 232386 584960 232476
rect 580441 232384 584960 232386
rect 580441 232328 580446 232384
rect 580502 232328 584960 232384
rect 580441 232326 584960 232328
rect 580441 232323 580507 232326
rect 583520 232236 584960 232326
rect 583520 218908 584960 219148
rect 583520 205580 584960 205820
rect 97717 196890 97783 196893
rect 99422 196890 100004 196924
rect 97717 196888 100004 196890
rect 97717 196832 97722 196888
rect 97778 196864 100004 196888
rect 97778 196832 99482 196864
rect 97717 196830 99482 196832
rect 97717 196827 97783 196830
rect 297265 196890 297331 196893
rect 299430 196890 300012 196924
rect 297265 196888 300012 196890
rect 297265 196832 297270 196888
rect 297326 196864 300012 196888
rect 297326 196832 299490 196864
rect 297265 196830 299490 196832
rect 297265 196827 297331 196830
rect 299054 196012 299060 196076
rect 299124 196074 299130 196076
rect 299381 196074 299447 196077
rect 299124 196072 299447 196074
rect 299124 196016 299386 196072
rect 299442 196016 299447 196072
rect 299124 196014 299447 196016
rect 299124 196012 299130 196014
rect 299381 196011 299447 196014
rect 97809 195938 97875 195941
rect 99422 195938 100004 195972
rect 97809 195936 100004 195938
rect 97809 195880 97814 195936
rect 97870 195912 100004 195936
rect 97870 195880 99482 195912
rect 97809 195878 99482 195880
rect 97809 195875 97875 195878
rect 297357 195938 297423 195941
rect 299614 195938 300012 195972
rect 297357 195936 300012 195938
rect 297357 195880 297362 195936
rect 297418 195912 300012 195936
rect 297418 195880 299674 195912
rect 297357 195878 299674 195880
rect 297357 195875 297423 195878
rect 294873 195258 294939 195261
rect 295190 195258 295196 195260
rect 294873 195256 295196 195258
rect 294873 195200 294878 195256
rect 294934 195200 295196 195256
rect 294873 195198 295196 195200
rect 294873 195195 294939 195198
rect 295190 195196 295196 195198
rect 295260 195196 295266 195260
rect 97809 193762 97875 193765
rect 99422 193762 100004 193796
rect 97809 193760 100004 193762
rect 97809 193704 97814 193760
rect 97870 193736 100004 193760
rect 97870 193704 99482 193736
rect 97809 193702 99482 193704
rect 97809 193699 97875 193702
rect 297449 193762 297515 193765
rect 299430 193762 300012 193796
rect 297449 193760 300012 193762
rect 297449 193704 297454 193760
rect 297510 193736 300012 193760
rect 297510 193704 299490 193736
rect 297449 193702 299490 193704
rect 297449 193699 297515 193702
rect 97717 192810 97783 192813
rect 99422 192810 100004 192844
rect 97717 192808 100004 192810
rect 97717 192752 97722 192808
rect 97778 192784 100004 192808
rect 97778 192752 99482 192784
rect 97717 192750 99482 192752
rect 97717 192747 97783 192750
rect 299013 192810 299079 192813
rect 299430 192810 300012 192844
rect 299013 192808 300012 192810
rect 299013 192752 299018 192808
rect 299074 192784 300012 192808
rect 299074 192752 299490 192784
rect 299013 192750 299490 192752
rect 299013 192747 299079 192750
rect 580349 192538 580415 192541
rect 583520 192538 584960 192628
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect 97533 191042 97599 191045
rect 99422 191042 100004 191076
rect 97533 191040 100004 191042
rect 97533 190984 97538 191040
rect 97594 191016 100004 191040
rect 97594 190984 99482 191016
rect 97533 190982 99482 190984
rect 97533 190979 97599 190982
rect 297541 191042 297607 191045
rect 299430 191042 300012 191076
rect 297541 191040 300012 191042
rect 297541 190984 297546 191040
rect 297602 191016 300012 191040
rect 297602 190984 299490 191016
rect 297541 190982 299490 190984
rect 297541 190979 297607 190982
rect 97625 189954 97691 189957
rect 99422 189954 100004 189988
rect 97625 189952 100004 189954
rect 97625 189896 97630 189952
rect 97686 189928 100004 189952
rect 97686 189896 99482 189928
rect 97625 189894 99482 189896
rect 97625 189891 97691 189894
rect -960 188866 480 188956
rect 3141 188866 3207 188869
rect -960 188864 3207 188866
rect -960 188808 3146 188864
rect 3202 188808 3207 188864
rect -960 188806 3207 188808
rect -960 188716 480 188806
rect 3141 188803 3207 188806
rect 297633 189954 297699 189957
rect 299430 189954 300012 189988
rect 297633 189952 300012 189954
rect 297633 189896 297638 189952
rect 297694 189928 300012 189952
rect 297694 189896 299490 189928
rect 297633 189894 299490 189896
rect 297633 189891 297699 189894
rect 297357 189138 297423 189141
rect 297633 189138 297699 189141
rect 297357 189136 297699 189138
rect 297357 189080 297362 189136
rect 297418 189080 297638 189136
rect 297694 189080 297699 189136
rect 297357 189078 297699 189080
rect 297357 189075 297423 189078
rect 297633 189075 297699 189078
rect 97441 188186 97507 188189
rect 99422 188186 100004 188220
rect 97441 188184 100004 188186
rect 97441 188128 97446 188184
rect 97502 188160 100004 188184
rect 97502 188128 99482 188160
rect 97441 188126 99482 188128
rect 97441 188123 97507 188126
rect -960 175796 480 176036
rect 297541 188186 297607 188189
rect 299105 188186 299171 188189
rect 299430 188186 300012 188220
rect 297541 188184 300012 188186
rect 297541 188128 297546 188184
rect 297602 188128 299110 188184
rect 299166 188160 300012 188184
rect 299166 188128 299490 188160
rect 297541 188126 299490 188128
rect 297541 188123 297607 188126
rect 299105 188123 299171 188126
rect 240133 175946 240199 175949
rect 277158 175946 277164 175948
rect 240133 175944 277164 175946
rect 240133 175888 240138 175944
rect 240194 175888 277164 175944
rect 240133 175886 277164 175888
rect 240133 175883 240199 175886
rect 277158 175884 277164 175886
rect 277228 175884 277234 175948
rect 583520 179060 584960 179300
rect 97349 169962 97415 169965
rect 99422 169962 100004 169996
rect 97349 169960 100004 169962
rect 97349 169904 97354 169960
rect 97410 169936 100004 169960
rect 97410 169904 99482 169936
rect 97349 169902 99482 169904
rect 97349 169899 97415 169902
rect 97901 168466 97967 168469
rect 97766 168464 97967 168466
rect 97766 168408 97906 168464
rect 97962 168408 97967 168464
rect 97766 168406 97967 168408
rect 97766 168194 97826 168406
rect 97901 168403 97967 168406
rect 297633 169962 297699 169965
rect 299430 169962 300012 169996
rect 297633 169960 300012 169962
rect 297633 169904 297638 169960
rect 297694 169936 300012 169960
rect 297694 169904 299490 169936
rect 297633 169902 299490 169904
rect 297633 169899 297699 169902
rect 97901 168330 97967 168333
rect 99422 168330 100004 168364
rect 97901 168328 100004 168330
rect 97901 168272 97906 168328
rect 97962 168304 100004 168328
rect 97962 168272 99482 168304
rect 97901 168270 99482 168272
rect 97901 168267 97967 168270
rect 97766 168134 99482 168194
rect 99422 168092 99482 168134
rect 297909 168330 297975 168333
rect 299430 168330 300012 168364
rect 297909 168328 300012 168330
rect 297909 168272 297914 168328
rect 297970 168304 300012 168328
rect 297970 168272 299490 168304
rect 297909 168270 299490 168272
rect 297909 168267 297975 168270
rect 99422 168032 100004 168092
rect -960 162890 480 162980
rect 3509 162890 3575 162893
rect -960 162888 3575 162890
rect -960 162832 3514 162888
rect 3570 162832 3575 162888
rect -960 162830 3575 162832
rect -960 162740 480 162830
rect 3509 162827 3575 162830
rect 297725 168058 297791 168061
rect 299430 168058 300012 168092
rect 297725 168056 300012 168058
rect 297725 168000 297730 168056
rect 297786 168032 300012 168056
rect 297786 168000 299490 168032
rect 297725 167998 299490 168000
rect 297725 167995 297791 167998
rect 293534 167044 293540 167108
rect 293604 167106 293610 167108
rect 293769 167106 293835 167109
rect 293604 167104 293835 167106
rect 293604 167048 293774 167104
rect 293830 167048 293835 167104
rect 293604 167046 293835 167048
rect 293604 167044 293610 167046
rect 293769 167043 293835 167046
rect 583520 165732 584960 165972
rect 158529 159900 158595 159901
rect 165981 159900 166047 159901
rect 158480 159898 158486 159900
rect 158438 159838 158486 159898
rect 158550 159896 158595 159900
rect 165960 159898 165966 159900
rect 158590 159840 158595 159896
rect 158480 159836 158486 159838
rect 158550 159836 158595 159840
rect 165890 159838 165966 159898
rect 166030 159896 166047 159900
rect 166042 159840 166047 159896
rect 165960 159836 165966 159838
rect 166030 159836 166047 159840
rect 158529 159835 158595 159836
rect 165981 159835 166047 159836
rect 173433 159900 173499 159901
rect 173433 159896 173446 159900
rect 173510 159898 173516 159900
rect 288985 159898 289051 159901
rect 316125 159898 316191 159901
rect 173433 159840 173438 159896
rect 173433 159836 173446 159840
rect 173510 159838 173590 159898
rect 288985 159896 316191 159898
rect 288985 159840 288990 159896
rect 289046 159840 316130 159896
rect 316186 159840 316191 159896
rect 288985 159838 316191 159840
rect 173510 159836 173516 159838
rect 173433 159835 173499 159836
rect 288985 159835 289051 159838
rect 316125 159835 316191 159838
rect 335997 159900 336063 159901
rect 338481 159900 338547 159901
rect 348233 159900 348299 159901
rect 335997 159896 336046 159900
rect 336110 159898 336116 159900
rect 335997 159840 336002 159896
rect 335997 159836 336046 159840
rect 336110 159838 336154 159898
rect 338481 159896 338494 159900
rect 338558 159898 338564 159900
rect 338481 159840 338486 159896
rect 336110 159836 336116 159838
rect 338481 159836 338494 159840
rect 338558 159838 338638 159898
rect 348233 159896 348286 159900
rect 348350 159898 348356 159900
rect 351913 159898 351979 159901
rect 348233 159840 348238 159896
rect 338558 159836 338564 159838
rect 348233 159836 348286 159840
rect 348350 159838 348390 159898
rect 348558 159896 351979 159898
rect 348558 159840 351918 159896
rect 351974 159840 351979 159896
rect 348558 159838 351979 159840
rect 348350 159836 348356 159838
rect 335997 159835 336063 159836
rect 338481 159835 338547 159836
rect 348233 159835 348299 159836
rect 294321 159762 294387 159765
rect 348558 159762 348618 159838
rect 351913 159835 351979 159838
rect 363505 159900 363571 159901
rect 370957 159900 371023 159901
rect 363505 159896 363518 159900
rect 363582 159898 363588 159900
rect 363505 159840 363510 159896
rect 363505 159836 363518 159840
rect 363582 159838 363662 159898
rect 370957 159896 370998 159900
rect 371062 159898 371068 159900
rect 370957 159840 370962 159896
rect 363582 159836 363588 159838
rect 370957 159836 370998 159840
rect 371062 159838 371114 159898
rect 371062 159836 371068 159838
rect 363505 159835 363571 159836
rect 370957 159835 371023 159836
rect 294321 159760 348618 159762
rect 294321 159704 294326 159760
rect 294382 159704 348618 159760
rect 294321 159702 348618 159704
rect 350993 159764 351059 159765
rect 353569 159764 353635 159765
rect 356053 159764 356119 159765
rect 360929 159764 360995 159765
rect 350993 159760 351006 159764
rect 351070 159762 351076 159764
rect 350993 159704 350998 159760
rect 294321 159699 294387 159702
rect 350993 159700 351006 159704
rect 351070 159702 351150 159762
rect 353569 159760 353590 159764
rect 353654 159762 353660 159764
rect 356032 159762 356038 159764
rect 353569 159704 353574 159760
rect 351070 159700 351076 159702
rect 353569 159700 353590 159704
rect 353654 159702 353726 159762
rect 355962 159702 356038 159762
rect 356102 159760 356119 159764
rect 356114 159704 356119 159760
rect 353654 159700 353660 159702
rect 356032 159700 356038 159702
rect 356102 159700 356119 159704
rect 360928 159700 360934 159764
rect 360998 159762 361004 159764
rect 360998 159702 361086 159762
rect 360998 159700 361004 159702
rect 350993 159699 351059 159700
rect 353569 159699 353635 159700
rect 356053 159699 356119 159700
rect 360929 159699 360995 159700
rect 156045 159628 156111 159629
rect 206001 159628 206067 159629
rect 156032 159626 156038 159628
rect 155954 159566 156038 159626
rect 156102 159624 156111 159628
rect 205944 159626 205950 159628
rect 156106 159568 156111 159624
rect 156032 159564 156038 159566
rect 156102 159564 156111 159568
rect 205910 159566 205950 159626
rect 206014 159624 206067 159628
rect 206062 159568 206067 159624
rect 205944 159564 205950 159566
rect 206014 159564 206067 159568
rect 156045 159563 156111 159564
rect 206001 159563 206067 159564
rect 298461 159626 298527 159629
rect 373993 159626 374059 159629
rect 298461 159624 374059 159626
rect 298461 159568 298466 159624
rect 298522 159568 373998 159624
rect 374054 159568 374059 159624
rect 298461 159566 374059 159568
rect 298461 159563 298527 159566
rect 373993 159563 374059 159566
rect 231853 159490 231919 159493
rect 275461 159490 275527 159493
rect 231853 159488 275527 159490
rect 231853 159432 231858 159488
rect 231914 159432 275466 159488
rect 275522 159432 275527 159488
rect 231853 159430 275527 159432
rect 231853 159427 231919 159430
rect 275461 159427 275527 159430
rect 298277 159490 298343 159493
rect 376753 159490 376819 159493
rect 298277 159488 376819 159490
rect 298277 159432 298282 159488
rect 298338 159432 376758 159488
rect 376814 159432 376819 159488
rect 298277 159430 376819 159432
rect 298277 159427 298343 159430
rect 376753 159427 376819 159430
rect 213913 159354 213979 159357
rect 273478 159354 273484 159356
rect 213913 159352 273484 159354
rect 213913 159296 213918 159352
rect 213974 159296 273484 159352
rect 213913 159294 273484 159296
rect 213913 159291 213979 159294
rect 273478 159292 273484 159294
rect 273548 159292 273554 159356
rect 298318 159292 298324 159356
rect 298388 159354 298394 159356
rect 378133 159354 378199 159357
rect 298388 159352 378199 159354
rect 298388 159296 378138 159352
rect 378194 159296 378199 159352
rect 298388 159294 378199 159296
rect 298388 159292 298394 159294
rect 378133 159291 378199 159294
rect 163630 159020 163636 159084
rect 163700 159082 163706 159084
rect 286174 159082 286180 159084
rect 163700 159022 286180 159082
rect 163700 159020 163706 159022
rect 286174 159020 286180 159022
rect 286244 159020 286250 159084
rect 153694 158884 153700 158948
rect 153764 158946 153770 158948
rect 283414 158946 283420 158948
rect 153764 158886 283420 158946
rect 153764 158884 153770 158886
rect 283414 158884 283420 158886
rect 283484 158884 283490 158948
rect 128302 158748 128308 158812
rect 128372 158810 128378 158812
rect 284702 158810 284708 158812
rect 128372 158750 284708 158810
rect 128372 158748 128378 158750
rect 284702 158748 284708 158750
rect 284772 158748 284778 158812
rect 286358 158748 286364 158812
rect 286428 158810 286434 158812
rect 286961 158810 287027 158813
rect 286428 158808 287027 158810
rect 286428 158752 286966 158808
rect 287022 158752 287027 158808
rect 286428 158750 287027 158752
rect 286428 158748 286434 158750
rect 286961 158747 287027 158750
rect 287646 158748 287652 158812
rect 287716 158810 287722 158812
rect 288341 158810 288407 158813
rect 287716 158808 288407 158810
rect 287716 158752 288346 158808
rect 288402 158752 288407 158808
rect 287716 158750 288407 158752
rect 287716 158748 287722 158750
rect 288341 158747 288407 158750
rect 288750 158748 288756 158812
rect 288820 158810 288826 158812
rect 289721 158810 289787 158813
rect 290641 158812 290707 158813
rect 290590 158810 290596 158812
rect 288820 158808 289787 158810
rect 288820 158752 289726 158808
rect 289782 158752 289787 158808
rect 288820 158750 289787 158752
rect 290550 158750 290596 158810
rect 290660 158808 290707 158812
rect 290702 158752 290707 158808
rect 288820 158748 288826 158750
rect 289721 158747 289787 158750
rect 290590 158748 290596 158750
rect 290660 158748 290707 158752
rect 290774 158748 290780 158812
rect 290844 158810 290850 158812
rect 291101 158810 291167 158813
rect 290844 158808 291167 158810
rect 290844 158752 291106 158808
rect 291162 158752 291167 158808
rect 290844 158750 291167 158752
rect 290844 158748 290850 158750
rect 290641 158747 290707 158748
rect 291101 158747 291167 158750
rect 291878 158748 291884 158812
rect 291948 158810 291954 158812
rect 292481 158810 292547 158813
rect 291948 158808 292547 158810
rect 291948 158752 292486 158808
rect 292542 158752 292547 158808
rect 291948 158750 292547 158752
rect 291948 158748 291954 158750
rect 292481 158747 292547 158750
rect 293350 158748 293356 158812
rect 293420 158810 293426 158812
rect 293493 158810 293559 158813
rect 295057 158812 295123 158813
rect 295006 158810 295012 158812
rect 293420 158808 293559 158810
rect 293420 158752 293498 158808
rect 293554 158752 293559 158808
rect 293420 158750 293559 158752
rect 294966 158750 295012 158810
rect 295076 158808 295123 158812
rect 295118 158752 295123 158808
rect 293420 158748 293426 158750
rect 293493 158747 293559 158750
rect 295006 158748 295012 158750
rect 295076 158748 295123 158752
rect 295926 158748 295932 158812
rect 295996 158810 296002 158812
rect 296621 158810 296687 158813
rect 295996 158808 296687 158810
rect 295996 158752 296626 158808
rect 296682 158752 296687 158808
rect 295996 158750 296687 158752
rect 295996 158748 296002 158750
rect 295057 158747 295123 158748
rect 296621 158747 296687 158750
rect 116158 158612 116164 158676
rect 116228 158674 116234 158676
rect 116485 158674 116551 158677
rect 116228 158672 116551 158674
rect 116228 158616 116490 158672
rect 116546 158616 116551 158672
rect 116228 158614 116551 158616
rect 116228 158612 116234 158614
rect 116485 158611 116551 158614
rect 117078 158612 117084 158676
rect 117148 158674 117154 158676
rect 117221 158674 117287 158677
rect 119705 158676 119771 158677
rect 120625 158676 120691 158677
rect 121913 158676 121979 158677
rect 123201 158676 123267 158677
rect 126513 158676 126579 158677
rect 119654 158674 119660 158676
rect 117148 158672 117287 158674
rect 117148 158616 117226 158672
rect 117282 158616 117287 158672
rect 117148 158614 117287 158616
rect 119614 158614 119660 158674
rect 119724 158672 119771 158676
rect 120574 158674 120580 158676
rect 119766 158616 119771 158672
rect 117148 158612 117154 158614
rect 117221 158611 117287 158614
rect 119654 158612 119660 158614
rect 119724 158612 119771 158616
rect 120534 158614 120580 158674
rect 120644 158672 120691 158676
rect 121862 158674 121868 158676
rect 120686 158616 120691 158672
rect 120574 158612 120580 158614
rect 120644 158612 120691 158616
rect 121822 158614 121868 158674
rect 121932 158672 121979 158676
rect 123150 158674 123156 158676
rect 121974 158616 121979 158672
rect 121862 158612 121868 158614
rect 121932 158612 121979 158616
rect 123110 158614 123156 158674
rect 123220 158672 123267 158676
rect 126462 158674 126468 158676
rect 123262 158616 123267 158672
rect 123150 158612 123156 158614
rect 123220 158612 123267 158616
rect 126422 158614 126468 158674
rect 126532 158672 126579 158676
rect 126574 158616 126579 158672
rect 126462 158612 126468 158614
rect 126532 158612 126579 158616
rect 127566 158612 127572 158676
rect 127636 158674 127642 158676
rect 128169 158674 128235 158677
rect 128721 158676 128787 158677
rect 128670 158674 128676 158676
rect 127636 158672 128235 158674
rect 127636 158616 128174 158672
rect 128230 158616 128235 158672
rect 127636 158614 128235 158616
rect 128630 158614 128676 158674
rect 128740 158672 128787 158676
rect 128782 158616 128787 158672
rect 127636 158612 127642 158614
rect 119705 158611 119771 158612
rect 120625 158611 120691 158612
rect 121913 158611 121979 158612
rect 123201 158611 123267 158612
rect 126513 158611 126579 158612
rect 128169 158611 128235 158614
rect 128670 158612 128676 158614
rect 128740 158612 128787 158616
rect 130142 158612 130148 158676
rect 130212 158674 130218 158676
rect 130561 158674 130627 158677
rect 130212 158672 130627 158674
rect 130212 158616 130566 158672
rect 130622 158616 130627 158672
rect 130212 158614 130627 158616
rect 130212 158612 130218 158614
rect 128721 158611 128787 158612
rect 130561 158611 130627 158614
rect 131246 158612 131252 158676
rect 131316 158674 131322 158676
rect 131481 158674 131547 158677
rect 132401 158676 132467 158677
rect 133505 158676 133571 158677
rect 132350 158674 132356 158676
rect 131316 158672 131547 158674
rect 131316 158616 131486 158672
rect 131542 158616 131547 158672
rect 131316 158614 131547 158616
rect 132310 158614 132356 158674
rect 132420 158672 132467 158676
rect 133454 158674 133460 158676
rect 132462 158616 132467 158672
rect 131316 158612 131322 158614
rect 131481 158611 131547 158614
rect 132350 158612 132356 158614
rect 132420 158612 132467 158616
rect 133414 158614 133460 158674
rect 133524 158672 133571 158676
rect 133566 158616 133571 158672
rect 133454 158612 133460 158614
rect 133524 158612 133571 158616
rect 134558 158612 134564 158676
rect 134628 158674 134634 158676
rect 134885 158674 134951 158677
rect 134628 158672 134951 158674
rect 134628 158616 134890 158672
rect 134946 158616 134951 158672
rect 134628 158614 134951 158616
rect 134628 158612 134634 158614
rect 132401 158611 132467 158612
rect 133505 158611 133571 158612
rect 134885 158611 134951 158614
rect 158110 158612 158116 158676
rect 158180 158674 158186 158676
rect 158529 158674 158595 158677
rect 158180 158672 158595 158674
rect 158180 158616 158534 158672
rect 158590 158616 158595 158672
rect 158180 158614 158595 158616
rect 158180 158612 158186 158614
rect 158529 158611 158595 158614
rect 159214 158612 159220 158676
rect 159284 158674 159290 158676
rect 159909 158674 159975 158677
rect 160921 158676 160987 158677
rect 168281 158676 168347 158677
rect 160870 158674 160876 158676
rect 159284 158672 159975 158674
rect 159284 158616 159914 158672
rect 159970 158616 159975 158672
rect 159284 158614 159975 158616
rect 160830 158614 160876 158674
rect 160940 158672 160987 158676
rect 168230 158674 168236 158676
rect 160982 158616 160987 158672
rect 159284 158612 159290 158614
rect 159909 158611 159975 158614
rect 160870 158612 160876 158614
rect 160940 158612 160987 158616
rect 168190 158614 168236 158674
rect 168300 158672 168347 158676
rect 168342 158616 168347 158672
rect 168230 158612 168236 158614
rect 168300 158612 168347 158616
rect 160921 158611 160987 158612
rect 168281 158611 168347 158612
rect 277945 158674 278011 158677
rect 278630 158674 278636 158676
rect 277945 158672 278636 158674
rect 277945 158616 277950 158672
rect 278006 158616 278636 158672
rect 277945 158614 278636 158616
rect 277945 158611 278011 158614
rect 278630 158612 278636 158614
rect 278700 158612 278706 158676
rect 315798 158612 315804 158676
rect 315868 158674 315874 158676
rect 316033 158674 316099 158677
rect 315868 158672 316099 158674
rect 315868 158616 316038 158672
rect 316094 158616 316099 158672
rect 315868 158614 316099 158616
rect 315868 158612 315874 158614
rect 316033 158611 316099 158614
rect 316953 158674 317019 158677
rect 318149 158676 318215 158677
rect 319437 158676 319503 158677
rect 320541 158676 320607 158677
rect 321645 158676 321711 158677
rect 323117 158676 323183 158677
rect 326429 158676 326495 158677
rect 328269 158676 328335 158677
rect 329925 158676 329991 158677
rect 317086 158674 317092 158676
rect 316953 158672 317092 158674
rect 316953 158616 316958 158672
rect 317014 158616 317092 158672
rect 316953 158614 317092 158616
rect 316953 158611 317019 158614
rect 317086 158612 317092 158614
rect 317156 158612 317162 158676
rect 318149 158672 318196 158676
rect 318260 158674 318266 158676
rect 318149 158616 318154 158672
rect 318149 158612 318196 158616
rect 318260 158614 318306 158674
rect 319437 158672 319484 158676
rect 319548 158674 319554 158676
rect 319437 158616 319442 158672
rect 318260 158612 318266 158614
rect 319437 158612 319484 158616
rect 319548 158614 319594 158674
rect 320541 158672 320588 158676
rect 320652 158674 320658 158676
rect 320541 158616 320546 158672
rect 319548 158612 319554 158614
rect 320541 158612 320588 158616
rect 320652 158614 320698 158674
rect 321645 158672 321692 158676
rect 321756 158674 321762 158676
rect 321645 158616 321650 158672
rect 320652 158612 320658 158614
rect 321645 158612 321692 158616
rect 321756 158614 321802 158674
rect 323117 158672 323164 158676
rect 323228 158674 323234 158676
rect 323117 158616 323122 158672
rect 321756 158612 321762 158614
rect 323117 158612 323164 158616
rect 323228 158614 323274 158674
rect 326429 158672 326476 158676
rect 326540 158674 326546 158676
rect 326429 158616 326434 158672
rect 323228 158612 323234 158614
rect 326429 158612 326476 158616
rect 326540 158614 326586 158674
rect 328269 158672 328316 158676
rect 328380 158674 328386 158676
rect 328269 158616 328274 158672
rect 326540 158612 326546 158614
rect 328269 158612 328316 158616
rect 328380 158614 328426 158674
rect 329925 158672 329972 158676
rect 330036 158674 330042 158676
rect 330569 158674 330635 158677
rect 333421 158676 333487 158677
rect 334525 158676 334591 158677
rect 330702 158674 330708 158676
rect 329925 158616 329930 158672
rect 328380 158612 328386 158614
rect 329925 158612 329972 158616
rect 330036 158614 330082 158674
rect 330569 158672 330708 158674
rect 330569 158616 330574 158672
rect 330630 158616 330708 158672
rect 330569 158614 330708 158616
rect 330036 158612 330042 158614
rect 318149 158611 318215 158612
rect 319437 158611 319503 158612
rect 320541 158611 320607 158612
rect 321645 158611 321711 158612
rect 323117 158611 323183 158612
rect 326429 158611 326495 158612
rect 328269 158611 328335 158612
rect 329925 158611 329991 158612
rect 330569 158611 330635 158614
rect 330702 158612 330708 158614
rect 330772 158612 330778 158676
rect 333421 158672 333468 158676
rect 333532 158674 333538 158676
rect 333421 158616 333426 158672
rect 333421 158612 333468 158616
rect 333532 158614 333578 158674
rect 334525 158672 334572 158676
rect 334636 158674 334642 158676
rect 335629 158674 335695 158677
rect 338113 158676 338179 158677
rect 335854 158674 335860 158676
rect 334525 158616 334530 158672
rect 333532 158612 333538 158614
rect 334525 158612 334572 158616
rect 334636 158614 334682 158674
rect 335629 158672 335860 158674
rect 335629 158616 335634 158672
rect 335690 158616 335860 158672
rect 335629 158614 335860 158616
rect 334636 158612 334642 158614
rect 333421 158611 333487 158612
rect 334525 158611 334591 158612
rect 335629 158611 335695 158614
rect 335854 158612 335860 158614
rect 335924 158612 335930 158676
rect 338062 158674 338068 158676
rect 338022 158614 338068 158674
rect 338132 158672 338179 158676
rect 338174 158616 338179 158672
rect 338062 158612 338068 158614
rect 338132 158612 338179 158616
rect 338113 158611 338179 158612
rect 340965 158676 341031 158677
rect 343541 158676 343607 158677
rect 343909 158676 343975 158677
rect 345933 158676 345999 158677
rect 348693 158676 348759 158677
rect 340965 158672 341012 158676
rect 341076 158674 341082 158676
rect 340965 158616 340970 158672
rect 340965 158612 341012 158616
rect 341076 158614 341122 158674
rect 343541 158672 343588 158676
rect 343652 158674 343658 158676
rect 343541 158616 343546 158672
rect 341076 158612 341082 158614
rect 343541 158612 343588 158616
rect 343652 158614 343698 158674
rect 343909 158672 343956 158676
rect 344020 158674 344026 158676
rect 343909 158616 343914 158672
rect 343652 158612 343658 158614
rect 343909 158612 343956 158616
rect 344020 158614 344066 158674
rect 345933 158672 345980 158676
rect 346044 158674 346050 158676
rect 345933 158616 345938 158672
rect 344020 158612 344026 158614
rect 345933 158612 345980 158616
rect 346044 158614 346090 158674
rect 348693 158672 348740 158676
rect 348804 158674 348810 158676
rect 355225 158674 355291 158677
rect 356973 158676 357039 158677
rect 358445 158676 358511 158677
rect 365805 158676 365871 158677
rect 368197 158676 368263 158677
rect 373349 158676 373415 158677
rect 376017 158676 376083 158677
rect 378593 158676 378659 158677
rect 380985 158676 381051 158677
rect 383561 158676 383627 158677
rect 385953 158676 386019 158677
rect 388529 158676 388595 158677
rect 355726 158674 355732 158676
rect 348693 158616 348698 158672
rect 346044 158612 346050 158614
rect 348693 158612 348740 158616
rect 348804 158614 348850 158674
rect 355225 158672 355732 158674
rect 355225 158616 355230 158672
rect 355286 158616 355732 158672
rect 355225 158614 355732 158616
rect 348804 158612 348810 158614
rect 340965 158611 341031 158612
rect 343541 158611 343607 158612
rect 343909 158611 343975 158612
rect 345933 158611 345999 158612
rect 348693 158611 348759 158612
rect 355225 158611 355291 158614
rect 355726 158612 355732 158614
rect 355796 158612 355802 158676
rect 356973 158672 357020 158676
rect 357084 158674 357090 158676
rect 356973 158616 356978 158672
rect 356973 158612 357020 158616
rect 357084 158614 357130 158674
rect 358445 158672 358492 158676
rect 358556 158674 358562 158676
rect 358445 158616 358450 158672
rect 357084 158612 357090 158614
rect 358445 158612 358492 158616
rect 358556 158614 358602 158674
rect 365805 158672 365852 158676
rect 365916 158674 365922 158676
rect 365805 158616 365810 158672
rect 358556 158612 358562 158614
rect 365805 158612 365852 158616
rect 365916 158614 365962 158674
rect 368197 158672 368244 158676
rect 368308 158674 368314 158676
rect 368197 158616 368202 158672
rect 365916 158612 365922 158614
rect 368197 158612 368244 158616
rect 368308 158614 368354 158674
rect 373349 158672 373396 158676
rect 373460 158674 373466 158676
rect 375966 158674 375972 158676
rect 373349 158616 373354 158672
rect 368308 158612 368314 158614
rect 373349 158612 373396 158616
rect 373460 158614 373506 158674
rect 375926 158614 375972 158674
rect 376036 158672 376083 158676
rect 378542 158674 378548 158676
rect 376078 158616 376083 158672
rect 373460 158612 373466 158614
rect 375966 158612 375972 158614
rect 376036 158612 376083 158616
rect 378502 158614 378548 158674
rect 378612 158672 378659 158676
rect 380934 158674 380940 158676
rect 378654 158616 378659 158672
rect 378542 158612 378548 158614
rect 378612 158612 378659 158616
rect 380894 158614 380940 158674
rect 381004 158672 381051 158676
rect 383510 158674 383516 158676
rect 381046 158616 381051 158672
rect 380934 158612 380940 158614
rect 381004 158612 381051 158616
rect 383470 158614 383516 158674
rect 383580 158672 383627 158676
rect 385902 158674 385908 158676
rect 383622 158616 383627 158672
rect 383510 158612 383516 158614
rect 383580 158612 383627 158616
rect 385862 158614 385908 158674
rect 385972 158672 386019 158676
rect 388478 158674 388484 158676
rect 386014 158616 386019 158672
rect 385902 158612 385908 158614
rect 385972 158612 386019 158616
rect 388438 158614 388484 158674
rect 388548 158672 388595 158676
rect 388590 158616 388595 158672
rect 388478 158612 388484 158614
rect 388548 158612 388595 158616
rect 391054 158612 391060 158676
rect 391124 158674 391130 158676
rect 391473 158674 391539 158677
rect 391124 158672 391539 158674
rect 391124 158616 391478 158672
rect 391534 158616 391539 158672
rect 391124 158614 391539 158616
rect 391124 158612 391130 158614
rect 356973 158611 357039 158612
rect 358445 158611 358511 158612
rect 365805 158611 365871 158612
rect 368197 158611 368263 158612
rect 373349 158611 373415 158612
rect 376017 158611 376083 158612
rect 378593 158611 378659 158612
rect 380985 158611 381051 158612
rect 383561 158611 383627 158612
rect 385953 158611 386019 158612
rect 388529 158611 388595 158612
rect 391473 158611 391539 158614
rect 393446 158612 393452 158676
rect 393516 158674 393522 158676
rect 394233 158674 394299 158677
rect 395889 158676 395955 158677
rect 398465 158676 398531 158677
rect 401041 158676 401107 158677
rect 395838 158674 395844 158676
rect 393516 158672 394299 158674
rect 393516 158616 394238 158672
rect 394294 158616 394299 158672
rect 393516 158614 394299 158616
rect 395798 158614 395844 158674
rect 395908 158672 395955 158676
rect 398414 158674 398420 158676
rect 395950 158616 395955 158672
rect 393516 158612 393522 158614
rect 394233 158611 394299 158614
rect 395838 158612 395844 158614
rect 395908 158612 395955 158616
rect 398374 158614 398420 158674
rect 398484 158672 398531 158676
rect 400990 158674 400996 158676
rect 398526 158616 398531 158672
rect 398414 158612 398420 158614
rect 398484 158612 398531 158616
rect 400950 158614 400996 158674
rect 401060 158672 401107 158676
rect 401102 158616 401107 158672
rect 400990 158612 400996 158614
rect 401060 158612 401107 158616
rect 403382 158612 403388 158676
rect 403452 158674 403458 158676
rect 403985 158674 404051 158677
rect 403452 158672 404051 158674
rect 403452 158616 403990 158672
rect 404046 158616 404051 158672
rect 403452 158614 404051 158616
rect 403452 158612 403458 158614
rect 395889 158611 395955 158612
rect 398465 158611 398531 158612
rect 401041 158611 401107 158612
rect 403985 158611 404051 158614
rect 405958 158612 405964 158676
rect 406028 158674 406034 158676
rect 406469 158674 406535 158677
rect 406028 158672 406535 158674
rect 406028 158616 406474 158672
rect 406530 158616 406535 158672
rect 406028 158614 406535 158616
rect 406028 158612 406034 158614
rect 406469 158611 406535 158614
rect 135897 158540 135963 158541
rect 137001 158540 137067 158541
rect 138105 158540 138171 158541
rect 135846 158538 135852 158540
rect 135806 158478 135852 158538
rect 135916 158536 135963 158540
rect 136950 158538 136956 158540
rect 135958 158480 135963 158536
rect 135846 158476 135852 158478
rect 135916 158476 135963 158480
rect 136910 158478 136956 158538
rect 137020 158536 137067 158540
rect 138054 158538 138060 158540
rect 137062 158480 137067 158536
rect 136950 158476 136956 158478
rect 137020 158476 137067 158480
rect 138014 158478 138060 158538
rect 138124 158536 138171 158540
rect 138166 158480 138171 158536
rect 138054 158476 138060 158478
rect 138124 158476 138171 158480
rect 148726 158476 148732 158540
rect 148796 158538 148802 158540
rect 148869 158538 148935 158541
rect 195881 158540 195947 158541
rect 195830 158538 195836 158540
rect 148796 158536 148935 158538
rect 148796 158480 148874 158536
rect 148930 158480 148935 158536
rect 148796 158478 148935 158480
rect 195790 158478 195836 158538
rect 195900 158536 195947 158540
rect 195942 158480 195947 158536
rect 148796 158476 148802 158478
rect 135897 158475 135963 158476
rect 137001 158475 137067 158476
rect 138105 158475 138171 158476
rect 148869 158475 148935 158478
rect 195830 158476 195836 158478
rect 195900 158476 195947 158480
rect 195881 158475 195947 158476
rect 276013 158538 276079 158541
rect 277025 158538 277091 158541
rect 358118 158538 358124 158540
rect 276013 158536 358124 158538
rect 276013 158480 276018 158536
rect 276074 158480 277030 158536
rect 277086 158480 358124 158536
rect 276013 158478 358124 158480
rect 276013 158475 276079 158478
rect 277025 158475 277091 158478
rect 358118 158476 358124 158478
rect 358188 158476 358194 158540
rect 118233 158404 118299 158405
rect 118182 158402 118188 158404
rect 118142 158342 118188 158402
rect 118252 158400 118299 158404
rect 118294 158344 118299 158400
rect 118182 158340 118188 158342
rect 118252 158340 118299 158344
rect 178534 158340 178540 158404
rect 178604 158402 178610 158404
rect 178861 158402 178927 158405
rect 178604 158400 178927 158402
rect 178604 158344 178866 158400
rect 178922 158344 178927 158400
rect 178604 158342 178927 158344
rect 178604 158340 178610 158342
rect 118233 158339 118299 158340
rect 178861 158339 178927 158342
rect 180926 158340 180932 158404
rect 180996 158402 181002 158404
rect 181805 158402 181871 158405
rect 180996 158400 181871 158402
rect 180996 158344 181810 158400
rect 181866 158344 181871 158400
rect 180996 158342 181871 158344
rect 180996 158340 181002 158342
rect 181805 158339 181871 158342
rect 183502 158340 183508 158404
rect 183572 158402 183578 158404
rect 184013 158402 184079 158405
rect 183572 158400 184079 158402
rect 183572 158344 184018 158400
rect 184074 158344 184079 158400
rect 183572 158342 184079 158344
rect 183572 158340 183578 158342
rect 184013 158339 184079 158342
rect 191046 158340 191052 158404
rect 191116 158402 191122 158404
rect 269849 158402 269915 158405
rect 191116 158400 269915 158402
rect 191116 158344 269854 158400
rect 269910 158344 269915 158400
rect 191116 158342 269915 158344
rect 191116 158340 191122 158342
rect 269849 158339 269915 158342
rect 271597 158402 271663 158405
rect 333605 158404 333671 158405
rect 332358 158402 332364 158404
rect 271597 158400 332364 158402
rect 271597 158344 271602 158400
rect 271658 158344 332364 158400
rect 271597 158342 332364 158344
rect 271597 158339 271663 158342
rect 332358 158340 332364 158342
rect 332428 158340 332434 158404
rect 333605 158400 333652 158404
rect 333716 158402 333722 158404
rect 336825 158402 336891 158405
rect 336958 158402 336964 158404
rect 333605 158344 333610 158400
rect 333605 158340 333652 158344
rect 333716 158342 333762 158402
rect 336825 158400 336964 158402
rect 336825 158344 336830 158400
rect 336886 158344 336964 158400
rect 336825 158342 336964 158344
rect 333716 158340 333722 158342
rect 333605 158339 333671 158340
rect 336825 158339 336891 158342
rect 336958 158340 336964 158342
rect 337028 158340 337034 158404
rect 141182 158204 141188 158268
rect 141252 158266 141258 158268
rect 141417 158266 141483 158269
rect 141785 158268 141851 158269
rect 141734 158266 141740 158268
rect 141252 158264 141483 158266
rect 141252 158208 141422 158264
rect 141478 158208 141483 158264
rect 141252 158206 141483 158208
rect 141694 158206 141740 158266
rect 141804 158264 141851 158268
rect 141846 158208 141851 158264
rect 141252 158204 141258 158206
rect 141417 158203 141483 158206
rect 141734 158204 141740 158206
rect 141804 158204 141851 158208
rect 143942 158204 143948 158268
rect 144012 158266 144018 158268
rect 144085 158266 144151 158269
rect 146017 158268 146083 158269
rect 146385 158268 146451 158269
rect 150985 158268 151051 158269
rect 185945 158268 186011 158269
rect 145966 158266 145972 158268
rect 144012 158264 144151 158266
rect 144012 158208 144090 158264
rect 144146 158208 144151 158264
rect 144012 158206 144151 158208
rect 145926 158206 145972 158266
rect 146036 158264 146083 158268
rect 146334 158266 146340 158268
rect 146078 158208 146083 158264
rect 144012 158204 144018 158206
rect 141785 158203 141851 158204
rect 144085 158203 144151 158206
rect 145966 158204 145972 158206
rect 146036 158204 146083 158208
rect 146294 158206 146340 158266
rect 146404 158264 146451 158268
rect 150934 158266 150940 158268
rect 146446 158208 146451 158264
rect 146334 158204 146340 158206
rect 146404 158204 146451 158208
rect 150894 158206 150940 158266
rect 151004 158264 151051 158268
rect 185894 158266 185900 158268
rect 151046 158208 151051 158264
rect 150934 158204 150940 158206
rect 151004 158204 151051 158208
rect 185854 158206 185900 158266
rect 185964 158264 186011 158268
rect 186006 158208 186011 158264
rect 185894 158204 185900 158206
rect 185964 158204 186011 158208
rect 193438 158204 193444 158268
rect 193508 158266 193514 158268
rect 270033 158266 270099 158269
rect 193508 158264 270099 158266
rect 193508 158208 270038 158264
rect 270094 158208 270099 158264
rect 193508 158206 270099 158208
rect 193508 158204 193514 158206
rect 146017 158203 146083 158204
rect 146385 158203 146451 158204
rect 150985 158203 151051 158204
rect 185945 158203 186011 158204
rect 270033 158203 270099 158206
rect 271689 158266 271755 158269
rect 331254 158266 331260 158268
rect 271689 158264 331260 158266
rect 271689 158208 271694 158264
rect 271750 158208 331260 158264
rect 271689 158206 331260 158208
rect 271689 158203 271755 158206
rect 331254 158204 331260 158206
rect 331324 158204 331330 158268
rect 338205 158266 338271 158269
rect 353293 158268 353359 158269
rect 339350 158266 339356 158268
rect 338205 158264 339356 158266
rect 338205 158208 338210 158264
rect 338266 158208 339356 158264
rect 338205 158206 339356 158208
rect 338205 158203 338271 158206
rect 339350 158204 339356 158206
rect 339420 158204 339426 158268
rect 353293 158264 353340 158268
rect 353404 158266 353410 158268
rect 353293 158208 353298 158264
rect 353293 158204 353340 158208
rect 353404 158206 353450 158266
rect 353404 158204 353410 158206
rect 353293 158203 353359 158204
rect 133689 158132 133755 158133
rect 133638 158130 133644 158132
rect 133598 158070 133644 158130
rect 133708 158128 133755 158132
rect 133750 158072 133755 158128
rect 133638 158068 133644 158070
rect 133708 158068 133755 158072
rect 170990 158068 170996 158132
rect 171060 158130 171066 158132
rect 238293 158130 238359 158133
rect 171060 158128 238359 158130
rect 171060 158072 238298 158128
rect 238354 158072 238359 158128
rect 171060 158070 238359 158072
rect 171060 158068 171066 158070
rect 133689 158067 133755 158068
rect 238293 158067 238359 158070
rect 274449 158130 274515 158133
rect 328678 158130 328684 158132
rect 274449 158128 328684 158130
rect 274449 158072 274454 158128
rect 274510 158072 328684 158128
rect 274449 158070 328684 158072
rect 274449 158067 274515 158070
rect 328678 158068 328684 158070
rect 328748 158068 328754 158132
rect 140681 157996 140747 157997
rect 140630 157994 140636 157996
rect 140590 157934 140636 157994
rect 140700 157992 140747 157996
rect 140742 157936 140747 157992
rect 140630 157932 140636 157934
rect 140700 157932 140747 157936
rect 188654 157932 188660 157996
rect 188724 157994 188730 157996
rect 238477 157994 238543 157997
rect 327574 157994 327580 157996
rect 188724 157992 238543 157994
rect 188724 157936 238482 157992
rect 238538 157936 238543 157992
rect 188724 157934 238543 157936
rect 188724 157932 188730 157934
rect 140681 157931 140747 157932
rect 238477 157931 238543 157934
rect 277350 157934 327580 157994
rect 136081 157860 136147 157861
rect 136030 157858 136036 157860
rect 135990 157798 136036 157858
rect 136100 157856 136147 157860
rect 136142 157800 136147 157856
rect 136030 157796 136036 157798
rect 136100 157796 136147 157800
rect 139526 157796 139532 157860
rect 139596 157858 139602 157860
rect 140497 157858 140563 157861
rect 145281 157860 145347 157861
rect 147673 157860 147739 157861
rect 145230 157858 145236 157860
rect 139596 157856 140563 157858
rect 139596 157800 140502 157856
rect 140558 157800 140563 157856
rect 139596 157798 140563 157800
rect 145190 157798 145236 157858
rect 145300 157856 145347 157860
rect 147622 157858 147628 157860
rect 145342 157800 145347 157856
rect 139596 157796 139602 157798
rect 136081 157795 136147 157796
rect 140497 157795 140563 157798
rect 145230 157796 145236 157798
rect 145300 157796 145347 157800
rect 147582 157798 147628 157858
rect 147692 157856 147739 157860
rect 147734 157800 147739 157856
rect 147622 157796 147628 157798
rect 147692 157796 147739 157800
rect 145281 157795 145347 157796
rect 147673 157795 147739 157796
rect 274357 157858 274423 157861
rect 277350 157858 277410 157934
rect 327574 157932 327580 157934
rect 327644 157932 327650 157996
rect 339493 157994 339559 157997
rect 340638 157994 340644 157996
rect 339493 157992 340644 157994
rect 339493 157936 339498 157992
rect 339554 157936 340644 157992
rect 339493 157934 340644 157936
rect 339493 157931 339559 157934
rect 340638 157932 340644 157934
rect 340708 157932 340714 157996
rect 342345 157994 342411 157997
rect 342846 157994 342852 157996
rect 342345 157992 342852 157994
rect 342345 157936 342350 157992
rect 342406 157936 342852 157992
rect 342345 157934 342852 157936
rect 342345 157931 342411 157934
rect 342846 157932 342852 157934
rect 342916 157932 342922 157996
rect 346669 157994 346735 157997
rect 347630 157994 347636 157996
rect 346669 157992 347636 157994
rect 346669 157936 346674 157992
rect 346730 157936 347636 157992
rect 346669 157934 347636 157936
rect 346669 157931 346735 157934
rect 347630 157932 347636 157934
rect 347700 157932 347706 157996
rect 274357 157856 277410 157858
rect 274357 157800 274362 157856
rect 274418 157800 277410 157856
rect 274357 157798 277410 157800
rect 324221 157860 324287 157861
rect 324221 157856 324268 157860
rect 324332 157858 324338 157860
rect 341057 157858 341123 157861
rect 341742 157858 341748 157860
rect 324221 157800 324226 157856
rect 274357 157795 274423 157798
rect 324221 157796 324268 157800
rect 324332 157798 324378 157858
rect 341057 157856 341748 157858
rect 341057 157800 341062 157856
rect 341118 157800 341748 157856
rect 341057 157798 341748 157800
rect 324332 157796 324338 157798
rect 324221 157795 324287 157796
rect 341057 157795 341123 157798
rect 341742 157796 341748 157798
rect 341812 157796 341818 157860
rect 345105 157858 345171 157861
rect 346393 157860 346459 157861
rect 345238 157858 345244 157860
rect 345105 157856 345244 157858
rect 345105 157800 345110 157856
rect 345166 157800 345244 157856
rect 345105 157798 345244 157800
rect 345105 157795 345171 157798
rect 345238 157796 345244 157798
rect 345308 157796 345314 157860
rect 346342 157858 346348 157860
rect 346302 157798 346348 157858
rect 346412 157856 346459 157860
rect 346454 157800 346459 157856
rect 346342 157796 346348 157798
rect 346412 157796 346459 157800
rect 346393 157795 346459 157796
rect 130694 157660 130700 157724
rect 130764 157722 130770 157724
rect 271413 157722 271479 157725
rect 130764 157720 271479 157722
rect 130764 157664 271418 157720
rect 271474 157664 271479 157720
rect 130764 157662 271479 157664
rect 130764 157660 130770 157662
rect 271413 157659 271479 157662
rect 124254 157524 124260 157588
rect 124324 157586 124330 157588
rect 124581 157586 124647 157589
rect 124324 157584 124647 157586
rect 124324 157528 124586 157584
rect 124642 157528 124647 157584
rect 124324 157526 124647 157528
rect 124324 157524 124330 157526
rect 124581 157523 124647 157526
rect 142838 157524 142844 157588
rect 142908 157586 142914 157588
rect 143073 157586 143139 157589
rect 198457 157588 198523 157589
rect 201033 157588 201099 157589
rect 203425 157588 203491 157589
rect 198406 157586 198412 157588
rect 142908 157584 143139 157586
rect 142908 157528 143078 157584
rect 143134 157528 143139 157584
rect 142908 157526 143139 157528
rect 198366 157526 198412 157586
rect 198476 157584 198523 157588
rect 200982 157586 200988 157588
rect 198518 157528 198523 157584
rect 142908 157524 142914 157526
rect 143073 157523 143139 157526
rect 198406 157524 198412 157526
rect 198476 157524 198523 157528
rect 200942 157526 200988 157586
rect 201052 157584 201099 157588
rect 203374 157586 203380 157588
rect 201094 157528 201099 157584
rect 200982 157524 200988 157526
rect 201052 157524 201099 157528
rect 203334 157526 203380 157586
rect 203444 157584 203491 157588
rect 203486 157528 203491 157584
rect 203374 157524 203380 157526
rect 203444 157524 203491 157528
rect 198457 157523 198523 157524
rect 201033 157523 201099 157524
rect 203425 157523 203491 157524
rect 274633 157586 274699 157589
rect 275921 157586 275987 157589
rect 359222 157586 359228 157588
rect 274633 157584 359228 157586
rect 274633 157528 274638 157584
rect 274694 157528 275926 157584
rect 275982 157528 359228 157584
rect 274633 157526 359228 157528
rect 274633 157523 274699 157526
rect 275921 157523 275987 157526
rect 359222 157524 359228 157526
rect 359292 157524 359298 157588
rect 125409 157452 125475 157453
rect 125358 157450 125364 157452
rect 125318 157390 125364 157450
rect 125428 157448 125475 157452
rect 125470 157392 125475 157448
rect 125358 157388 125364 157390
rect 125428 157388 125475 157392
rect 138606 157388 138612 157452
rect 138676 157388 138682 157452
rect 143574 157388 143580 157452
rect 143644 157450 143650 157452
rect 144361 157450 144427 157453
rect 143644 157448 144427 157450
rect 143644 157392 144366 157448
rect 144422 157392 144427 157448
rect 143644 157390 144427 157392
rect 143644 157388 143650 157390
rect 125409 157387 125475 157388
rect 138614 157314 138674 157388
rect 144361 157387 144427 157390
rect 148358 157388 148364 157452
rect 148428 157450 148434 157452
rect 148501 157450 148567 157453
rect 149881 157452 149947 157453
rect 151353 157452 151419 157453
rect 149830 157450 149836 157452
rect 148428 157448 148567 157450
rect 148428 157392 148506 157448
rect 148562 157392 148567 157448
rect 148428 157390 148567 157392
rect 149790 157390 149836 157450
rect 149900 157448 149947 157452
rect 151302 157450 151308 157452
rect 149942 157392 149947 157448
rect 148428 157388 148434 157390
rect 148501 157387 148567 157390
rect 149830 157388 149836 157390
rect 149900 157388 149947 157392
rect 151262 157390 151308 157450
rect 151372 157448 151419 157452
rect 151414 157392 151419 157448
rect 151302 157388 151308 157390
rect 151372 157388 151419 157392
rect 152222 157388 152228 157452
rect 152292 157450 152298 157452
rect 152641 157450 152707 157453
rect 152292 157448 152707 157450
rect 152292 157392 152646 157448
rect 152702 157392 152707 157448
rect 152292 157390 152707 157392
rect 152292 157388 152298 157390
rect 149881 157387 149947 157388
rect 151353 157387 151419 157388
rect 152641 157387 152707 157390
rect 153326 157388 153332 157452
rect 153396 157450 153402 157452
rect 154113 157450 154179 157453
rect 154481 157452 154547 157453
rect 155769 157452 155835 157453
rect 157057 157452 157123 157453
rect 154430 157450 154436 157452
rect 153396 157448 154179 157450
rect 153396 157392 154118 157448
rect 154174 157392 154179 157448
rect 153396 157390 154179 157392
rect 154390 157390 154436 157450
rect 154500 157448 154547 157452
rect 155718 157450 155724 157452
rect 154542 157392 154547 157448
rect 153396 157388 153402 157390
rect 154113 157387 154179 157390
rect 154430 157388 154436 157390
rect 154500 157388 154547 157392
rect 155678 157390 155724 157450
rect 155788 157448 155835 157452
rect 157006 157450 157012 157452
rect 155830 157392 155835 157448
rect 155718 157388 155724 157390
rect 155788 157388 155835 157392
rect 156966 157390 157012 157450
rect 157076 157448 157123 157452
rect 157118 157392 157123 157448
rect 157006 157388 157012 157390
rect 157076 157388 157123 157392
rect 175958 157388 175964 157452
rect 176028 157450 176034 157452
rect 280889 157450 280955 157453
rect 176028 157448 280955 157450
rect 176028 157392 280894 157448
rect 280950 157392 280955 157448
rect 176028 157390 280955 157392
rect 176028 157388 176034 157390
rect 154481 157387 154547 157388
rect 155769 157387 155835 157388
rect 157057 157387 157123 157388
rect 280889 157387 280955 157390
rect 291694 157388 291700 157452
rect 291764 157450 291770 157452
rect 292389 157450 292455 157453
rect 291764 157448 292455 157450
rect 291764 157392 292394 157448
rect 292450 157392 292455 157448
rect 291764 157390 292455 157392
rect 291764 157388 291770 157390
rect 292389 157387 292455 157390
rect 325325 157452 325391 157453
rect 349797 157452 349863 157453
rect 325325 157448 325372 157452
rect 325436 157450 325442 157452
rect 325325 157392 325330 157448
rect 325325 157388 325372 157392
rect 325436 157390 325482 157450
rect 349797 157448 349844 157452
rect 349908 157450 349914 157452
rect 350993 157450 351059 157453
rect 352189 157452 352255 157453
rect 354397 157452 354463 157453
rect 351126 157450 351132 157452
rect 349797 157392 349802 157448
rect 325436 157388 325442 157390
rect 349797 157388 349844 157392
rect 349908 157390 349954 157450
rect 350993 157448 351132 157450
rect 350993 157392 350998 157448
rect 351054 157392 351132 157448
rect 350993 157390 351132 157392
rect 349908 157388 349914 157390
rect 325325 157387 325391 157388
rect 349797 157387 349863 157388
rect 350993 157387 351059 157390
rect 351126 157388 351132 157390
rect 351196 157388 351202 157452
rect 352189 157448 352236 157452
rect 352300 157450 352306 157452
rect 352189 157392 352194 157448
rect 352189 157388 352236 157392
rect 352300 157390 352346 157450
rect 354397 157448 354444 157452
rect 354508 157450 354514 157452
rect 354397 157392 354402 157448
rect 352300 157388 352306 157390
rect 354397 157388 354444 157392
rect 354508 157390 354554 157450
rect 354508 157388 354514 157390
rect 352189 157387 352255 157388
rect 354397 157387 354463 157388
rect 261661 157314 261727 157317
rect 138614 157312 261727 157314
rect 138614 157256 261666 157312
rect 261722 157256 261727 157312
rect 138614 157254 261727 157256
rect 261661 157251 261727 157254
rect 202873 156906 202939 156909
rect 270953 156906 271019 156909
rect 202873 156904 271019 156906
rect 202873 156848 202878 156904
rect 202934 156848 270958 156904
rect 271014 156848 271019 156904
rect 202873 156846 271019 156848
rect 202873 156843 202939 156846
rect 270953 156843 271019 156846
rect 175273 156770 175339 156773
rect 256049 156770 256115 156773
rect 175273 156768 256115 156770
rect 175273 156712 175278 156768
rect 175334 156712 256054 156768
rect 256110 156712 256115 156768
rect 175273 156710 256115 156712
rect 175273 156707 175339 156710
rect 256049 156707 256115 156710
rect 144913 156634 144979 156637
rect 262673 156634 262739 156637
rect 144913 156632 262739 156634
rect 144913 156576 144918 156632
rect 144974 156576 262678 156632
rect 262734 156576 262739 156632
rect 144913 156574 262739 156576
rect 144913 156571 144979 156574
rect 262673 156571 262739 156574
rect 133689 155954 133755 155957
rect 264421 155954 264487 155957
rect 133689 155952 264487 155954
rect 133689 155896 133694 155952
rect 133750 155896 264426 155952
rect 264482 155896 264487 155952
rect 133689 155894 264487 155896
rect 133689 155891 133755 155894
rect 264421 155891 264487 155894
rect 220813 155546 220879 155549
rect 273621 155546 273687 155549
rect 220813 155544 273687 155546
rect 220813 155488 220818 155544
rect 220874 155488 273626 155544
rect 273682 155488 273687 155544
rect 220813 155486 273687 155488
rect 220813 155483 220879 155486
rect 273621 155483 273687 155486
rect 178033 155410 178099 155413
rect 268285 155410 268351 155413
rect 178033 155408 268351 155410
rect 178033 155352 178038 155408
rect 178094 155352 268290 155408
rect 268346 155352 268351 155408
rect 178033 155350 268351 155352
rect 178033 155347 178099 155350
rect 268285 155347 268351 155350
rect 153193 155274 153259 155277
rect 257429 155274 257495 155277
rect 153193 155272 257495 155274
rect 153193 155216 153198 155272
rect 153254 155216 257434 155272
rect 257490 155216 257495 155272
rect 153193 155214 257495 155216
rect 153193 155211 153259 155214
rect 257429 155211 257495 155214
rect 287830 155212 287836 155276
rect 287900 155274 287906 155276
rect 309133 155274 309199 155277
rect 287900 155272 309199 155274
rect 287900 155216 309138 155272
rect 309194 155216 309199 155272
rect 287900 155214 309199 155216
rect 287900 155212 287906 155214
rect 309133 155211 309199 155214
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect 195973 152418 196039 152421
rect 270534 152418 270540 152420
rect 195973 152416 270540 152418
rect 195973 152360 195978 152416
rect 196034 152360 270540 152416
rect 195973 152358 270540 152360
rect 195973 152355 196039 152358
rect 270534 152356 270540 152358
rect 270604 152356 270610 152420
rect 298134 152356 298140 152420
rect 298204 152418 298210 152420
rect 380893 152418 380959 152421
rect 298204 152416 380959 152418
rect 298204 152360 380898 152416
rect 380954 152360 380959 152416
rect 298204 152358 380959 152360
rect 298204 152356 298210 152358
rect 380893 152355 380959 152358
rect 268469 151058 268535 151061
rect 278814 151058 278820 151060
rect 268469 151056 278820 151058
rect 268469 151000 268474 151056
rect 268530 151000 278820 151056
rect 268469 150998 278820 151000
rect 268469 150995 268535 150998
rect 278814 150996 278820 150998
rect 278884 150996 278890 151060
rect -960 149834 480 149924
rect 3601 149834 3667 149837
rect -960 149832 3667 149834
rect -960 149776 3606 149832
rect 3662 149776 3667 149832
rect -960 149774 3667 149776
rect -960 149684 480 149774
rect 3601 149771 3667 149774
rect 293166 149092 293172 149156
rect 293236 149154 293242 149156
rect 293585 149154 293651 149157
rect 293236 149152 293651 149154
rect 293236 149096 293590 149152
rect 293646 149096 293651 149152
rect 293236 149094 293651 149096
rect 293236 149092 293242 149094
rect 293585 149091 293651 149094
rect 293718 148276 293724 148340
rect 293788 148338 293794 148340
rect 345013 148338 345079 148341
rect 293788 148336 345079 148338
rect 293788 148280 345018 148336
rect 345074 148280 345079 148336
rect 293788 148278 345079 148280
rect 293788 148276 293794 148278
rect 345013 148275 345079 148278
rect 222193 146978 222259 146981
rect 274766 146978 274772 146980
rect 222193 146976 274772 146978
rect 222193 146920 222198 146976
rect 222254 146920 274772 146976
rect 222193 146918 274772 146920
rect 222193 146915 222259 146918
rect 274766 146916 274772 146918
rect 274836 146916 274842 146980
rect 583520 139212 584960 139452
rect 215293 138682 215359 138685
rect 273294 138682 273300 138684
rect 215293 138680 273300 138682
rect 215293 138624 215298 138680
rect 215354 138624 273300 138680
rect 215293 138622 273300 138624
rect 215293 138619 215359 138622
rect 273294 138620 273300 138622
rect 273364 138620 273370 138684
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 223573 127666 223639 127669
rect 274582 127666 274588 127668
rect 223573 127664 274588 127666
rect 223573 127608 223578 127664
rect 223634 127608 274588 127664
rect 223573 127606 274588 127608
rect 223573 127603 223639 127606
rect 274582 127604 274588 127606
rect 274652 127604 274658 127668
rect 583520 125884 584960 126124
rect 282177 125490 282243 125493
rect 282862 125490 282868 125492
rect 282177 125488 282868 125490
rect 282177 125432 282182 125488
rect 282238 125432 282868 125488
rect 282177 125430 282868 125432
rect 282177 125427 282243 125430
rect 282862 125428 282868 125430
rect 282932 125428 282938 125492
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 298502 82044 298508 82108
rect 298572 82106 298578 82108
rect 379513 82106 379579 82109
rect 298572 82104 379579 82106
rect 298572 82048 379518 82104
rect 379574 82048 379579 82104
rect 298572 82046 379579 82048
rect 298572 82044 298578 82046
rect 379513 82043 379579 82046
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 439446 71844 439452 71908
rect 439516 71906 439522 71908
rect 583526 71906 583586 72798
rect 439516 71846 583586 71906
rect 439516 71844 439522 71846
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect 282310 9556 282316 9620
rect 282380 9618 282386 9620
rect 364609 9618 364675 9621
rect 282380 9616 364675 9618
rect 282380 9560 364614 9616
rect 364670 9560 364675 9616
rect 282380 9558 364675 9560
rect 282380 9556 282386 9558
rect 364609 9555 364675 9558
rect 279918 9420 279924 9484
rect 279988 9482 279994 9484
rect 370589 9482 370655 9485
rect 279988 9480 370655 9482
rect 279988 9424 370594 9480
rect 370650 9424 370655 9480
rect 279988 9422 370655 9424
rect 279988 9420 279994 9422
rect 370589 9419 370655 9422
rect 292246 9284 292252 9348
rect 292316 9346 292322 9348
rect 394233 9346 394299 9349
rect 292316 9344 394299 9346
rect 292316 9288 394238 9344
rect 394294 9288 394299 9344
rect 292316 9286 394299 9288
rect 292316 9284 292322 9286
rect 394233 9283 394299 9286
rect 283966 9148 283972 9212
rect 284036 9210 284042 9212
rect 401317 9210 401383 9213
rect 284036 9208 401383 9210
rect 284036 9152 401322 9208
rect 401378 9152 401383 9208
rect 284036 9150 401383 9152
rect 284036 9148 284042 9150
rect 401317 9147 401383 9150
rect 284886 9012 284892 9076
rect 284956 9074 284962 9076
rect 404813 9074 404879 9077
rect 284956 9072 404879 9074
rect 284956 9016 404818 9072
rect 404874 9016 404879 9072
rect 284956 9014 404879 9016
rect 284956 9012 284962 9014
rect 404813 9011 404879 9014
rect 284150 8876 284156 8940
rect 284220 8938 284226 8940
rect 411897 8938 411963 8941
rect 284220 8936 411963 8938
rect 284220 8880 411902 8936
rect 411958 8880 411963 8936
rect 284220 8878 411963 8880
rect 284220 8876 284226 8878
rect 411897 8875 411963 8878
rect 292430 8740 292436 8804
rect 292500 8802 292506 8804
rect 337469 8802 337535 8805
rect 292500 8800 337535 8802
rect 292500 8744 337474 8800
rect 337530 8744 337535 8800
rect 292500 8742 337535 8744
rect 292500 8740 292506 8742
rect 337469 8739 337535 8742
rect 296294 7516 296300 7580
rect 296364 7578 296370 7580
rect 362309 7578 362375 7581
rect 296364 7576 362375 7578
rect 296364 7520 362314 7576
rect 362370 7520 362375 7576
rect 296364 7518 362375 7520
rect 296364 7516 296370 7518
rect 362309 7515 362375 7518
rect 297766 6836 297772 6900
rect 297836 6898 297842 6900
rect 372889 6898 372955 6901
rect 297836 6896 372955 6898
rect 297836 6840 372894 6896
rect 372950 6840 372955 6896
rect 297836 6838 372955 6840
rect 297836 6836 297842 6838
rect 372889 6835 372955 6838
rect 289302 6700 289308 6764
rect 289372 6762 289378 6764
rect 382365 6762 382431 6765
rect 289372 6760 382431 6762
rect 289372 6704 382370 6760
rect 382426 6704 382431 6760
rect 289372 6702 382431 6704
rect 289372 6700 289378 6702
rect 382365 6699 382431 6702
rect -960 6490 480 6580
rect 289118 6564 289124 6628
rect 289188 6626 289194 6628
rect 385953 6626 386019 6629
rect 289188 6624 386019 6626
rect 289188 6568 385958 6624
rect 386014 6568 386019 6624
rect 289188 6566 386019 6568
rect 289188 6564 289194 6566
rect 385953 6563 386019 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 289486 6428 289492 6492
rect 289556 6490 289562 6492
rect 389449 6490 389515 6493
rect 289556 6488 389515 6490
rect 289556 6432 389454 6488
rect 389510 6432 389515 6488
rect 583520 6476 584960 6716
rect 289556 6430 389515 6432
rect 289556 6428 289562 6430
rect 389449 6427 389515 6430
rect 286726 6292 286732 6356
rect 286796 6354 286802 6356
rect 393037 6354 393103 6357
rect 286796 6352 393103 6354
rect 286796 6296 393042 6352
rect 393098 6296 393103 6352
rect 286796 6294 393103 6296
rect 286796 6292 286802 6294
rect 393037 6291 393103 6294
rect 288014 6156 288020 6220
rect 288084 6218 288090 6220
rect 396533 6218 396599 6221
rect 288084 6216 396599 6218
rect 288084 6160 396538 6216
rect 396594 6160 396599 6216
rect 288084 6158 396599 6160
rect 288084 6156 288090 6158
rect 396533 6155 396599 6158
rect 297582 6020 297588 6084
rect 297652 6082 297658 6084
rect 371693 6082 371759 6085
rect 297652 6080 371759 6082
rect 297652 6024 371698 6080
rect 371754 6024 371759 6080
rect 297652 6022 371759 6024
rect 297652 6020 297658 6022
rect 371693 6019 371759 6022
rect 296478 4932 296484 4996
rect 296548 4994 296554 4996
rect 363505 4994 363571 4997
rect 296548 4992 363571 4994
rect 296548 4936 363510 4992
rect 363566 4936 363571 4992
rect 296548 4934 363571 4936
rect 296548 4932 296554 4934
rect 363505 4931 363571 4934
rect 297950 4796 297956 4860
rect 298020 4858 298026 4860
rect 368197 4858 368263 4861
rect 298020 4856 368263 4858
rect 298020 4800 368202 4856
rect 368258 4800 368263 4856
rect 298020 4798 368263 4800
rect 298020 4796 298026 4798
rect 368197 4795 368263 4798
rect 282494 3980 282500 4044
rect 282564 4042 282570 4044
rect 356329 4042 356395 4045
rect 282564 4040 356395 4042
rect 282564 3984 356334 4040
rect 356390 3984 356395 4040
rect 282564 3982 356395 3984
rect 282564 3980 282570 3982
rect 356329 3979 356395 3982
rect 280470 3844 280476 3908
rect 280540 3906 280546 3908
rect 367001 3906 367067 3909
rect 280540 3904 367067 3906
rect 280540 3848 367006 3904
rect 367062 3848 367067 3904
rect 280540 3846 367067 3848
rect 280540 3844 280546 3846
rect 367001 3843 367067 3846
rect 296110 3708 296116 3772
rect 296180 3770 296186 3772
rect 388253 3770 388319 3773
rect 296180 3768 388319 3770
rect 296180 3712 388258 3768
rect 388314 3712 388319 3768
rect 296180 3710 388319 3712
rect 296180 3708 296186 3710
rect 388253 3707 388319 3710
rect 433241 3770 433307 3773
rect 440417 3770 440483 3773
rect 433241 3768 440483 3770
rect 433241 3712 433246 3768
rect 433302 3712 440422 3768
rect 440478 3712 440483 3768
rect 433241 3710 440483 3712
rect 433241 3707 433307 3710
rect 440417 3707 440483 3710
rect 286910 3572 286916 3636
rect 286980 3634 286986 3636
rect 383561 3634 383627 3637
rect 286980 3632 383627 3634
rect 286980 3576 383566 3632
rect 383622 3576 383627 3632
rect 286980 3574 383627 3576
rect 286980 3572 286986 3574
rect 383561 3571 383627 3574
rect 437422 3572 437428 3636
rect 437492 3634 437498 3636
rect 437933 3634 437999 3637
rect 437492 3632 437999 3634
rect 437492 3576 437938 3632
rect 437994 3576 437999 3632
rect 437492 3574 437999 3576
rect 437492 3572 437498 3574
rect 437933 3571 437999 3574
rect 288198 3436 288204 3500
rect 288268 3498 288274 3500
rect 387149 3498 387215 3501
rect 288268 3496 387215 3498
rect 288268 3440 387154 3496
rect 387210 3440 387215 3496
rect 288268 3438 387215 3440
rect 288268 3436 288274 3438
rect 387149 3435 387215 3438
rect 435541 3498 435607 3501
rect 439129 3500 439195 3501
rect 437606 3498 437612 3500
rect 435541 3496 437612 3498
rect 435541 3440 435546 3496
rect 435602 3440 437612 3496
rect 435541 3438 437612 3440
rect 435541 3435 435607 3438
rect 437606 3436 437612 3438
rect 437676 3436 437682 3500
rect 439078 3436 439084 3500
rect 439148 3498 439195 3500
rect 439148 3496 439240 3498
rect 439190 3440 439240 3496
rect 439148 3438 439240 3440
rect 439148 3436 439195 3438
rect 439129 3435 439195 3436
rect 258257 3362 258323 3365
rect 280286 3362 280292 3364
rect 258257 3360 280292 3362
rect 258257 3304 258262 3360
rect 258318 3304 280292 3360
rect 258257 3302 280292 3304
rect 258257 3299 258323 3302
rect 280286 3300 280292 3302
rect 280356 3300 280362 3364
rect 285070 3300 285076 3364
rect 285140 3362 285146 3364
rect 390645 3362 390711 3365
rect 285140 3360 390711 3362
rect 285140 3304 390650 3360
rect 390706 3304 390711 3360
rect 285140 3302 390711 3304
rect 285140 3300 285146 3302
rect 390645 3299 390711 3302
rect 434437 3362 434503 3365
rect 437790 3362 437796 3364
rect 434437 3360 437796 3362
rect 434437 3304 434442 3360
rect 434498 3304 437796 3360
rect 434437 3302 437796 3304
rect 434437 3299 434503 3302
rect 437790 3300 437796 3302
rect 437860 3300 437866 3364
rect 282678 3164 282684 3228
rect 282748 3226 282754 3228
rect 320909 3226 320975 3229
rect 282748 3224 320975 3226
rect 282748 3168 320914 3224
rect 320970 3168 320975 3224
rect 282748 3166 320975 3168
rect 282748 3164 282754 3166
rect 320909 3163 320975 3166
<< obsm3 >>
rect 220000 516924 356620 563308
rect 220064 516864 356620 516924
rect 220000 515972 356620 516864
rect 220064 515912 356620 515972
rect 220000 513796 356620 515912
rect 220064 513736 356620 513796
rect 220000 512844 356620 513736
rect 220064 512784 356620 512844
rect 220000 511076 356620 512784
rect 220064 511016 356620 511076
rect 220000 509988 356620 511016
rect 220064 509928 356620 509988
rect 220000 508220 356620 509928
rect 220064 508160 356620 508220
rect 220000 489996 356620 508160
rect 220064 489936 356620 489996
rect 220000 488364 356620 489936
rect 220064 488304 356620 488364
rect 220000 488092 356620 488304
rect 220064 488032 356620 488092
rect 220000 480000 356620 488032
rect 100000 196924 236620 243308
rect 300000 196924 436620 243308
rect 100004 196864 236620 196924
rect 100000 195972 236620 196864
rect 300012 196864 436620 196924
rect 300000 195972 436620 196864
rect 100004 195912 236620 195972
rect 100000 193796 236620 195912
rect 300012 195912 436620 195972
rect 300000 193796 436620 195912
rect 100004 193736 236620 193796
rect 100000 192844 236620 193736
rect 300012 193736 436620 193796
rect 300000 192844 436620 193736
rect 100004 192784 236620 192844
rect 100000 191076 236620 192784
rect 300012 192784 436620 192844
rect 300000 191076 436620 192784
rect 100004 191016 236620 191076
rect 100000 189988 236620 191016
rect 300012 191016 436620 191076
rect 300000 189988 436620 191016
rect 100004 189928 236620 189988
rect 100000 188220 236620 189928
rect 300012 189928 436620 189988
rect 300000 188220 436620 189928
rect 100004 188160 236620 188220
rect 100000 169996 236620 188160
rect 300012 188160 436620 188220
rect 300000 169996 436620 188160
rect 100004 169936 236620 169996
rect 100000 168364 236620 169936
rect 300012 169936 436620 169996
rect 300000 168364 436620 169936
rect 100004 168304 236620 168364
rect 100000 168092 236620 168304
rect 300012 168304 436620 168364
rect 300000 168092 436620 168304
rect 100004 168032 236620 168092
rect 100000 160000 236620 168032
rect 300012 168032 436620 168092
rect 300000 160000 436620 168032
<< via3 >>
rect 243124 477260 243188 477324
rect 254532 476988 254596 477052
rect 265940 476988 266004 477052
rect 270908 476988 270972 477052
rect 305868 476988 305932 477052
rect 308444 476988 308508 477052
rect 256188 476852 256252 476916
rect 278452 476852 278516 476916
rect 311020 476852 311084 476916
rect 323348 476852 323412 476916
rect 260972 476716 261036 476780
rect 303476 476716 303540 476780
rect 244228 476640 244292 476644
rect 244228 476584 244278 476640
rect 244278 476584 244292 476640
rect 244228 476580 244292 476584
rect 248276 476580 248340 476644
rect 253612 476580 253676 476644
rect 257844 476580 257908 476644
rect 258396 476580 258460 476644
rect 263548 476640 263612 476644
rect 263548 476584 263598 476640
rect 263598 476584 263612 476640
rect 263548 476580 263612 476584
rect 276060 476640 276124 476644
rect 276060 476584 276074 476640
rect 276074 476584 276124 476640
rect 276060 476580 276124 476584
rect 250668 476444 250732 476508
rect 268332 476444 268396 476508
rect 273484 476444 273548 476508
rect 313412 476444 313476 476508
rect 315804 476444 315868 476508
rect 237236 476368 237300 476372
rect 237236 476312 237286 476368
rect 237286 476312 237300 476368
rect 237236 476308 237300 476312
rect 245332 476308 245396 476372
rect 251404 476308 251468 476372
rect 260604 476308 260668 476372
rect 266492 476308 266556 476372
rect 273300 476308 273364 476372
rect 318380 476308 318444 476372
rect 320956 476308 321020 476372
rect 235948 476232 236012 476236
rect 235948 476176 235962 476232
rect 235962 476176 236012 476232
rect 235948 476172 236012 476176
rect 238156 476172 238220 476236
rect 239628 476172 239692 476236
rect 240548 476172 240612 476236
rect 241836 476172 241900 476236
rect 246436 476172 246500 476236
rect 247540 476172 247604 476236
rect 248644 476172 248708 476236
rect 250116 476172 250180 476236
rect 252324 476172 252388 476236
rect 253428 476172 253492 476236
rect 255820 476172 255884 476236
rect 257108 476172 257172 476236
rect 259500 476172 259564 476236
rect 261708 476172 261772 476236
rect 262812 476172 262876 476236
rect 263916 476172 263980 476236
rect 265388 476172 265452 476236
rect 267596 476232 267660 476236
rect 267596 476176 267610 476232
rect 267610 476176 267660 476232
rect 267596 476172 267660 476176
rect 268700 476172 268764 476236
rect 269804 476172 269868 476236
rect 271276 476172 271340 476236
rect 272196 476172 272260 476236
rect 274404 476172 274468 476236
rect 275876 476232 275940 476236
rect 275876 476176 275926 476232
rect 275926 476176 275940 476232
rect 275876 476172 275940 476176
rect 276980 476172 277044 476236
rect 278084 476172 278148 476236
rect 279188 476172 279252 476236
rect 280844 476172 280908 476236
rect 283420 476172 283484 476236
rect 285996 476172 286060 476236
rect 288204 476172 288268 476236
rect 290964 476172 291028 476236
rect 293356 476172 293420 476236
rect 295932 476172 295996 476236
rect 298508 476172 298572 476236
rect 300900 476232 300964 476236
rect 300900 476176 300914 476232
rect 300914 476176 300964 476232
rect 300900 476172 300964 476176
rect 325924 476172 325988 476236
rect 439452 444348 439516 444412
rect 286180 308756 286244 308820
rect 292436 308680 292500 308684
rect 292436 308624 292486 308680
rect 292486 308624 292500 308680
rect 292436 308620 292500 308624
rect 297956 308620 298020 308684
rect 270540 308272 270604 308276
rect 270540 308216 270590 308272
rect 270590 308216 270604 308272
rect 270540 308212 270604 308216
rect 284708 308212 284772 308276
rect 297772 308076 297836 308140
rect 298324 308076 298388 308140
rect 273300 307940 273364 308004
rect 274588 307940 274652 308004
rect 283420 307940 283484 308004
rect 273484 307804 273548 307868
rect 274772 307804 274836 307868
rect 277348 307864 277412 307868
rect 277348 307808 277398 307864
rect 277398 307808 277412 307864
rect 277348 307804 277412 307808
rect 278820 307864 278884 307868
rect 278820 307808 278870 307864
rect 278870 307808 278884 307864
rect 278820 307804 278884 307808
rect 280292 307804 280356 307868
rect 283052 307864 283116 307868
rect 283052 307808 283102 307864
rect 283102 307808 283116 307864
rect 283052 307804 283116 307808
rect 287836 307804 287900 307868
rect 293724 307864 293788 307868
rect 293724 307808 293774 307864
rect 293774 307808 293788 307864
rect 293724 307804 293788 307808
rect 296300 307864 296364 307868
rect 296300 307808 296350 307864
rect 296350 307808 296364 307864
rect 296300 307804 296364 307808
rect 296484 307864 296548 307868
rect 296484 307808 296534 307864
rect 296534 307808 296548 307864
rect 296484 307804 296548 307808
rect 297588 307804 297652 307868
rect 298508 307804 298572 307868
rect 278636 306172 278700 306236
rect 437428 297332 437492 297396
rect 439084 261428 439148 261492
rect 288204 248236 288268 248300
rect 437612 248236 437676 248300
rect 286916 248100 286980 248164
rect 282316 247964 282380 248028
rect 285076 247828 285140 247892
rect 279924 247692 279988 247756
rect 283972 247556 284036 247620
rect 292252 247420 292316 247484
rect 284156 247012 284220 247076
rect 284892 247012 284956 247076
rect 286364 247012 286428 247076
rect 287652 247012 287716 247076
rect 288756 247012 288820 247076
rect 293172 247012 293236 247076
rect 295012 247072 295076 247076
rect 295012 247016 295062 247072
rect 295062 247016 295076 247072
rect 295012 247012 295076 247016
rect 289308 245516 289372 245580
rect 289124 245380 289188 245444
rect 293540 245244 293604 245308
rect 298140 245516 298204 245580
rect 296116 245380 296180 245444
rect 437796 245244 437860 245308
rect 286732 245108 286796 245172
rect 282500 244972 282564 245036
rect 299060 245108 299124 245172
rect 280476 244836 280540 244900
rect 295196 244896 295260 244900
rect 295196 244840 295246 244896
rect 295246 244840 295260 244896
rect 295196 244836 295260 244840
rect 282684 244700 282748 244764
rect 293356 244760 293420 244764
rect 293356 244704 293406 244760
rect 293406 244704 293420 244760
rect 293356 244700 293420 244704
rect 295932 244700 295996 244764
rect 289492 244564 289556 244628
rect 290780 244488 290844 244492
rect 290780 244432 290830 244488
rect 290830 244432 290844 244488
rect 290780 244428 290844 244432
rect 288020 244292 288084 244356
rect 290596 244292 290660 244356
rect 291700 244352 291764 244356
rect 291700 244296 291750 244352
rect 291750 244296 291764 244352
rect 291700 244292 291764 244296
rect 291884 244292 291948 244356
rect 299060 196012 299124 196076
rect 295196 195196 295260 195260
rect 277164 175884 277228 175948
rect 293540 167044 293604 167108
rect 158486 159896 158550 159900
rect 158486 159840 158534 159896
rect 158534 159840 158550 159896
rect 158486 159836 158550 159840
rect 165966 159896 166030 159900
rect 165966 159840 165986 159896
rect 165986 159840 166030 159896
rect 165966 159836 166030 159840
rect 173446 159896 173510 159900
rect 173446 159840 173494 159896
rect 173494 159840 173510 159896
rect 173446 159836 173510 159840
rect 336046 159896 336110 159900
rect 336046 159840 336058 159896
rect 336058 159840 336110 159896
rect 336046 159836 336110 159840
rect 338494 159896 338558 159900
rect 338494 159840 338542 159896
rect 338542 159840 338558 159896
rect 338494 159836 338558 159840
rect 348286 159896 348350 159900
rect 348286 159840 348294 159896
rect 348294 159840 348350 159896
rect 348286 159836 348350 159840
rect 363518 159896 363582 159900
rect 363518 159840 363566 159896
rect 363566 159840 363582 159896
rect 363518 159836 363582 159840
rect 370998 159896 371062 159900
rect 370998 159840 371018 159896
rect 371018 159840 371062 159896
rect 370998 159836 371062 159840
rect 351006 159760 351070 159764
rect 351006 159704 351054 159760
rect 351054 159704 351070 159760
rect 351006 159700 351070 159704
rect 353590 159760 353654 159764
rect 353590 159704 353630 159760
rect 353630 159704 353654 159760
rect 353590 159700 353654 159704
rect 356038 159760 356102 159764
rect 356038 159704 356058 159760
rect 356058 159704 356102 159760
rect 356038 159700 356102 159704
rect 360934 159760 360998 159764
rect 360934 159704 360990 159760
rect 360990 159704 360998 159760
rect 360934 159700 360998 159704
rect 156038 159624 156102 159628
rect 156038 159568 156050 159624
rect 156050 159568 156102 159624
rect 156038 159564 156102 159568
rect 205950 159624 206014 159628
rect 205950 159568 206006 159624
rect 206006 159568 206014 159624
rect 205950 159564 206014 159568
rect 273484 159292 273548 159356
rect 298324 159292 298388 159356
rect 163636 159020 163700 159084
rect 286180 159020 286244 159084
rect 153700 158884 153764 158948
rect 283420 158884 283484 158948
rect 128308 158748 128372 158812
rect 284708 158748 284772 158812
rect 286364 158748 286428 158812
rect 287652 158748 287716 158812
rect 288756 158748 288820 158812
rect 290596 158808 290660 158812
rect 290596 158752 290646 158808
rect 290646 158752 290660 158808
rect 290596 158748 290660 158752
rect 290780 158748 290844 158812
rect 291884 158748 291948 158812
rect 293356 158748 293420 158812
rect 295012 158808 295076 158812
rect 295012 158752 295062 158808
rect 295062 158752 295076 158808
rect 295012 158748 295076 158752
rect 295932 158748 295996 158812
rect 116164 158612 116228 158676
rect 117084 158612 117148 158676
rect 119660 158672 119724 158676
rect 119660 158616 119710 158672
rect 119710 158616 119724 158672
rect 119660 158612 119724 158616
rect 120580 158672 120644 158676
rect 120580 158616 120630 158672
rect 120630 158616 120644 158672
rect 120580 158612 120644 158616
rect 121868 158672 121932 158676
rect 121868 158616 121918 158672
rect 121918 158616 121932 158672
rect 121868 158612 121932 158616
rect 123156 158672 123220 158676
rect 123156 158616 123206 158672
rect 123206 158616 123220 158672
rect 123156 158612 123220 158616
rect 126468 158672 126532 158676
rect 126468 158616 126518 158672
rect 126518 158616 126532 158672
rect 126468 158612 126532 158616
rect 127572 158612 127636 158676
rect 128676 158672 128740 158676
rect 128676 158616 128726 158672
rect 128726 158616 128740 158672
rect 128676 158612 128740 158616
rect 130148 158612 130212 158676
rect 131252 158612 131316 158676
rect 132356 158672 132420 158676
rect 132356 158616 132406 158672
rect 132406 158616 132420 158672
rect 132356 158612 132420 158616
rect 133460 158672 133524 158676
rect 133460 158616 133510 158672
rect 133510 158616 133524 158672
rect 133460 158612 133524 158616
rect 134564 158612 134628 158676
rect 158116 158612 158180 158676
rect 159220 158612 159284 158676
rect 160876 158672 160940 158676
rect 160876 158616 160926 158672
rect 160926 158616 160940 158672
rect 160876 158612 160940 158616
rect 168236 158672 168300 158676
rect 168236 158616 168286 158672
rect 168286 158616 168300 158672
rect 168236 158612 168300 158616
rect 278636 158612 278700 158676
rect 315804 158612 315868 158676
rect 317092 158612 317156 158676
rect 318196 158672 318260 158676
rect 318196 158616 318210 158672
rect 318210 158616 318260 158672
rect 318196 158612 318260 158616
rect 319484 158672 319548 158676
rect 319484 158616 319498 158672
rect 319498 158616 319548 158672
rect 319484 158612 319548 158616
rect 320588 158672 320652 158676
rect 320588 158616 320602 158672
rect 320602 158616 320652 158672
rect 320588 158612 320652 158616
rect 321692 158672 321756 158676
rect 321692 158616 321706 158672
rect 321706 158616 321756 158672
rect 321692 158612 321756 158616
rect 323164 158672 323228 158676
rect 323164 158616 323178 158672
rect 323178 158616 323228 158672
rect 323164 158612 323228 158616
rect 326476 158672 326540 158676
rect 326476 158616 326490 158672
rect 326490 158616 326540 158672
rect 326476 158612 326540 158616
rect 328316 158672 328380 158676
rect 328316 158616 328330 158672
rect 328330 158616 328380 158672
rect 328316 158612 328380 158616
rect 329972 158672 330036 158676
rect 329972 158616 329986 158672
rect 329986 158616 330036 158672
rect 329972 158612 330036 158616
rect 330708 158612 330772 158676
rect 333468 158672 333532 158676
rect 333468 158616 333482 158672
rect 333482 158616 333532 158672
rect 333468 158612 333532 158616
rect 334572 158672 334636 158676
rect 334572 158616 334586 158672
rect 334586 158616 334636 158672
rect 334572 158612 334636 158616
rect 335860 158612 335924 158676
rect 338068 158672 338132 158676
rect 338068 158616 338118 158672
rect 338118 158616 338132 158672
rect 338068 158612 338132 158616
rect 341012 158672 341076 158676
rect 341012 158616 341026 158672
rect 341026 158616 341076 158672
rect 341012 158612 341076 158616
rect 343588 158672 343652 158676
rect 343588 158616 343602 158672
rect 343602 158616 343652 158672
rect 343588 158612 343652 158616
rect 343956 158672 344020 158676
rect 343956 158616 343970 158672
rect 343970 158616 344020 158672
rect 343956 158612 344020 158616
rect 345980 158672 346044 158676
rect 345980 158616 345994 158672
rect 345994 158616 346044 158672
rect 345980 158612 346044 158616
rect 348740 158672 348804 158676
rect 348740 158616 348754 158672
rect 348754 158616 348804 158672
rect 348740 158612 348804 158616
rect 355732 158612 355796 158676
rect 357020 158672 357084 158676
rect 357020 158616 357034 158672
rect 357034 158616 357084 158672
rect 357020 158612 357084 158616
rect 358492 158672 358556 158676
rect 358492 158616 358506 158672
rect 358506 158616 358556 158672
rect 358492 158612 358556 158616
rect 365852 158672 365916 158676
rect 365852 158616 365866 158672
rect 365866 158616 365916 158672
rect 365852 158612 365916 158616
rect 368244 158672 368308 158676
rect 368244 158616 368258 158672
rect 368258 158616 368308 158672
rect 368244 158612 368308 158616
rect 373396 158672 373460 158676
rect 373396 158616 373410 158672
rect 373410 158616 373460 158672
rect 373396 158612 373460 158616
rect 375972 158672 376036 158676
rect 375972 158616 376022 158672
rect 376022 158616 376036 158672
rect 375972 158612 376036 158616
rect 378548 158672 378612 158676
rect 378548 158616 378598 158672
rect 378598 158616 378612 158672
rect 378548 158612 378612 158616
rect 380940 158672 381004 158676
rect 380940 158616 380990 158672
rect 380990 158616 381004 158672
rect 380940 158612 381004 158616
rect 383516 158672 383580 158676
rect 383516 158616 383566 158672
rect 383566 158616 383580 158672
rect 383516 158612 383580 158616
rect 385908 158672 385972 158676
rect 385908 158616 385958 158672
rect 385958 158616 385972 158672
rect 385908 158612 385972 158616
rect 388484 158672 388548 158676
rect 388484 158616 388534 158672
rect 388534 158616 388548 158672
rect 388484 158612 388548 158616
rect 391060 158612 391124 158676
rect 393452 158612 393516 158676
rect 395844 158672 395908 158676
rect 395844 158616 395894 158672
rect 395894 158616 395908 158672
rect 395844 158612 395908 158616
rect 398420 158672 398484 158676
rect 398420 158616 398470 158672
rect 398470 158616 398484 158672
rect 398420 158612 398484 158616
rect 400996 158672 401060 158676
rect 400996 158616 401046 158672
rect 401046 158616 401060 158672
rect 400996 158612 401060 158616
rect 403388 158612 403452 158676
rect 405964 158612 406028 158676
rect 135852 158536 135916 158540
rect 135852 158480 135902 158536
rect 135902 158480 135916 158536
rect 135852 158476 135916 158480
rect 136956 158536 137020 158540
rect 136956 158480 137006 158536
rect 137006 158480 137020 158536
rect 136956 158476 137020 158480
rect 138060 158536 138124 158540
rect 138060 158480 138110 158536
rect 138110 158480 138124 158536
rect 138060 158476 138124 158480
rect 148732 158476 148796 158540
rect 195836 158536 195900 158540
rect 195836 158480 195886 158536
rect 195886 158480 195900 158536
rect 195836 158476 195900 158480
rect 358124 158476 358188 158540
rect 118188 158400 118252 158404
rect 118188 158344 118238 158400
rect 118238 158344 118252 158400
rect 118188 158340 118252 158344
rect 178540 158340 178604 158404
rect 180932 158340 180996 158404
rect 183508 158340 183572 158404
rect 191052 158340 191116 158404
rect 332364 158340 332428 158404
rect 333652 158400 333716 158404
rect 333652 158344 333666 158400
rect 333666 158344 333716 158400
rect 333652 158340 333716 158344
rect 336964 158340 337028 158404
rect 141188 158204 141252 158268
rect 141740 158264 141804 158268
rect 141740 158208 141790 158264
rect 141790 158208 141804 158264
rect 141740 158204 141804 158208
rect 143948 158204 144012 158268
rect 145972 158264 146036 158268
rect 145972 158208 146022 158264
rect 146022 158208 146036 158264
rect 145972 158204 146036 158208
rect 146340 158264 146404 158268
rect 146340 158208 146390 158264
rect 146390 158208 146404 158264
rect 146340 158204 146404 158208
rect 150940 158264 151004 158268
rect 150940 158208 150990 158264
rect 150990 158208 151004 158264
rect 150940 158204 151004 158208
rect 185900 158264 185964 158268
rect 185900 158208 185950 158264
rect 185950 158208 185964 158264
rect 185900 158204 185964 158208
rect 193444 158204 193508 158268
rect 331260 158204 331324 158268
rect 339356 158204 339420 158268
rect 353340 158264 353404 158268
rect 353340 158208 353354 158264
rect 353354 158208 353404 158264
rect 353340 158204 353404 158208
rect 133644 158128 133708 158132
rect 133644 158072 133694 158128
rect 133694 158072 133708 158128
rect 133644 158068 133708 158072
rect 170996 158068 171060 158132
rect 328684 158068 328748 158132
rect 140636 157992 140700 157996
rect 140636 157936 140686 157992
rect 140686 157936 140700 157992
rect 140636 157932 140700 157936
rect 188660 157932 188724 157996
rect 136036 157856 136100 157860
rect 136036 157800 136086 157856
rect 136086 157800 136100 157856
rect 136036 157796 136100 157800
rect 139532 157796 139596 157860
rect 145236 157856 145300 157860
rect 145236 157800 145286 157856
rect 145286 157800 145300 157856
rect 145236 157796 145300 157800
rect 147628 157856 147692 157860
rect 147628 157800 147678 157856
rect 147678 157800 147692 157856
rect 147628 157796 147692 157800
rect 327580 157932 327644 157996
rect 340644 157932 340708 157996
rect 342852 157932 342916 157996
rect 347636 157932 347700 157996
rect 324268 157856 324332 157860
rect 324268 157800 324282 157856
rect 324282 157800 324332 157856
rect 324268 157796 324332 157800
rect 341748 157796 341812 157860
rect 345244 157796 345308 157860
rect 346348 157856 346412 157860
rect 346348 157800 346398 157856
rect 346398 157800 346412 157856
rect 346348 157796 346412 157800
rect 130700 157660 130764 157724
rect 124260 157524 124324 157588
rect 142844 157524 142908 157588
rect 198412 157584 198476 157588
rect 198412 157528 198462 157584
rect 198462 157528 198476 157584
rect 198412 157524 198476 157528
rect 200988 157584 201052 157588
rect 200988 157528 201038 157584
rect 201038 157528 201052 157584
rect 200988 157524 201052 157528
rect 203380 157584 203444 157588
rect 203380 157528 203430 157584
rect 203430 157528 203444 157584
rect 203380 157524 203444 157528
rect 359228 157524 359292 157588
rect 125364 157448 125428 157452
rect 125364 157392 125414 157448
rect 125414 157392 125428 157448
rect 125364 157388 125428 157392
rect 138612 157388 138676 157452
rect 143580 157388 143644 157452
rect 148364 157388 148428 157452
rect 149836 157448 149900 157452
rect 149836 157392 149886 157448
rect 149886 157392 149900 157448
rect 149836 157388 149900 157392
rect 151308 157448 151372 157452
rect 151308 157392 151358 157448
rect 151358 157392 151372 157448
rect 151308 157388 151372 157392
rect 152228 157388 152292 157452
rect 153332 157388 153396 157452
rect 154436 157448 154500 157452
rect 154436 157392 154486 157448
rect 154486 157392 154500 157448
rect 154436 157388 154500 157392
rect 155724 157448 155788 157452
rect 155724 157392 155774 157448
rect 155774 157392 155788 157448
rect 155724 157388 155788 157392
rect 157012 157448 157076 157452
rect 157012 157392 157062 157448
rect 157062 157392 157076 157448
rect 157012 157388 157076 157392
rect 175964 157388 176028 157452
rect 291700 157388 291764 157452
rect 325372 157448 325436 157452
rect 325372 157392 325386 157448
rect 325386 157392 325436 157448
rect 325372 157388 325436 157392
rect 349844 157448 349908 157452
rect 349844 157392 349858 157448
rect 349858 157392 349908 157448
rect 349844 157388 349908 157392
rect 351132 157388 351196 157452
rect 352236 157448 352300 157452
rect 352236 157392 352250 157448
rect 352250 157392 352300 157448
rect 352236 157388 352300 157392
rect 354444 157448 354508 157452
rect 354444 157392 354458 157448
rect 354458 157392 354508 157448
rect 354444 157388 354508 157392
rect 287836 155212 287900 155276
rect 270540 152356 270604 152420
rect 298140 152356 298204 152420
rect 278820 150996 278884 151060
rect 293172 149092 293236 149156
rect 293724 148276 293788 148340
rect 274772 146916 274836 146980
rect 273300 138620 273364 138684
rect 274588 127604 274652 127668
rect 282868 125428 282932 125492
rect 298508 82044 298572 82108
rect 439452 71844 439516 71908
rect 282316 9556 282380 9620
rect 279924 9420 279988 9484
rect 292252 9284 292316 9348
rect 283972 9148 284036 9212
rect 284892 9012 284956 9076
rect 284156 8876 284220 8940
rect 292436 8740 292500 8804
rect 296300 7516 296364 7580
rect 297772 6836 297836 6900
rect 289308 6700 289372 6764
rect 289124 6564 289188 6628
rect 289492 6428 289556 6492
rect 286732 6292 286796 6356
rect 288020 6156 288084 6220
rect 297588 6020 297652 6084
rect 296484 4932 296548 4996
rect 297956 4796 298020 4860
rect 282500 3980 282564 4044
rect 280476 3844 280540 3908
rect 296116 3708 296180 3772
rect 286916 3572 286980 3636
rect 437428 3572 437492 3636
rect 288204 3436 288268 3500
rect 437612 3436 437676 3500
rect 439084 3496 439148 3500
rect 439084 3440 439134 3496
rect 439134 3440 439148 3496
rect 439084 3436 439148 3440
rect 280292 3300 280356 3364
rect 285076 3300 285140 3364
rect 437796 3300 437860 3364
rect 282684 3164 282748 3228
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 245308 101414 245898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 245308 105914 250398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 245308 110414 254898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 245308 114914 259398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 245308 119414 263898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 245308 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 245308 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 245308 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 245308 137414 245898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 245308 141914 250398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 245308 146414 254898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 245308 150914 259398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 245308 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 245308 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 245308 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 245308 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 245308 173414 245898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 245308 177914 250398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 245308 182414 254898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 245308 186914 259398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 245308 191414 263898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 245308 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 245308 200414 272898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 245308 204914 277398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 245308 209414 245898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 565308 218414 578898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 565308 222914 583398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 565308 227414 587898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 565308 231914 592398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 565308 236414 596898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 565308 240914 565398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 565308 245414 569898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 565308 249914 574398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 565308 254414 578898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 565308 258914 583398
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 565308 263414 587898
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 565308 267914 592398
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 565308 272414 596898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 565308 276914 565398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 565308 281414 569898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 565308 285914 574398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 565308 290414 578898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 565308 294914 583398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 565308 299414 587898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 565308 303914 592398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 565308 308414 596898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 565308 312914 565398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 565308 317414 569898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 565308 321914 574398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 565308 326414 578898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 565308 330914 583398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 565308 335414 587898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 565308 339914 592398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 565308 344414 596898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 565308 348914 565398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 565308 353414 569898
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 565308 357914 574398
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 220272 547954 220620 547986
rect 220272 547718 220328 547954
rect 220564 547718 220620 547954
rect 220272 547634 220620 547718
rect 220272 547398 220328 547634
rect 220564 547398 220620 547634
rect 220272 547366 220620 547398
rect 356000 547954 356348 547986
rect 356000 547718 356056 547954
rect 356292 547718 356348 547954
rect 356000 547634 356348 547718
rect 356000 547398 356056 547634
rect 356292 547398 356348 547634
rect 356000 547366 356348 547398
rect 220952 543454 221300 543486
rect 220952 543218 221008 543454
rect 221244 543218 221300 543454
rect 220952 543134 221300 543218
rect 220952 542898 221008 543134
rect 221244 542898 221300 543134
rect 220952 542866 221300 542898
rect 355320 543454 355668 543486
rect 355320 543218 355376 543454
rect 355612 543218 355668 543454
rect 355320 543134 355668 543218
rect 355320 542898 355376 543134
rect 355612 542898 355668 543134
rect 355320 542866 355668 542898
rect 220272 511954 220620 511986
rect 220272 511718 220328 511954
rect 220564 511718 220620 511954
rect 220272 511634 220620 511718
rect 220272 511398 220328 511634
rect 220564 511398 220620 511634
rect 220272 511366 220620 511398
rect 356000 511954 356348 511986
rect 356000 511718 356056 511954
rect 356292 511718 356348 511954
rect 356000 511634 356348 511718
rect 356000 511398 356056 511634
rect 356292 511398 356348 511634
rect 356000 511366 356348 511398
rect 220952 507454 221300 507486
rect 220952 507218 221008 507454
rect 221244 507218 221300 507454
rect 220952 507134 221300 507218
rect 220952 506898 221008 507134
rect 221244 506898 221300 507134
rect 220952 506866 221300 506898
rect 355320 507454 355668 507486
rect 355320 507218 355376 507454
rect 355612 507218 355668 507454
rect 355320 507134 355668 507218
rect 355320 506898 355376 507134
rect 355612 506898 355668 507134
rect 355320 506866 355668 506898
rect 236056 479770 236116 480080
rect 235950 479710 236116 479770
rect 237144 479770 237204 480080
rect 238232 479770 238292 480080
rect 237144 479710 237298 479770
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 245308 213914 250398
rect 217794 471454 218414 478000
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 245308 218414 254898
rect 222294 475954 222914 478000
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 245308 222914 259398
rect 226794 444454 227414 478000
rect 235950 476237 236010 479710
rect 237238 476373 237298 479710
rect 238158 479710 238292 479770
rect 239592 479770 239652 480080
rect 240544 479770 240604 480080
rect 241768 479770 241828 480080
rect 243128 479770 243188 480080
rect 239592 479710 239690 479770
rect 240544 479710 240610 479770
rect 241768 479710 241898 479770
rect 237235 476372 237301 476373
rect 237235 476308 237236 476372
rect 237300 476308 237301 476372
rect 237235 476307 237301 476308
rect 238158 476237 238218 479710
rect 239630 476237 239690 479710
rect 240550 476237 240610 479710
rect 241838 476237 241898 479710
rect 243126 479710 243188 479770
rect 244216 479770 244276 480080
rect 245440 479770 245500 480080
rect 246528 479770 246588 480080
rect 247616 479770 247676 480080
rect 248296 479770 248356 480080
rect 248704 479770 248764 480080
rect 244216 479710 244290 479770
rect 243126 477325 243186 479710
rect 243123 477324 243189 477325
rect 243123 477260 243124 477324
rect 243188 477260 243189 477324
rect 243123 477259 243189 477260
rect 244230 476645 244290 479710
rect 245334 479710 245500 479770
rect 246438 479710 246588 479770
rect 247542 479710 247676 479770
rect 248278 479710 248356 479770
rect 248646 479710 248764 479770
rect 250064 479770 250124 480080
rect 250744 479770 250804 480080
rect 250064 479710 250178 479770
rect 244227 476644 244293 476645
rect 244227 476580 244228 476644
rect 244292 476580 244293 476644
rect 244227 476579 244293 476580
rect 245334 476373 245394 479710
rect 245331 476372 245397 476373
rect 245331 476308 245332 476372
rect 245396 476308 245397 476372
rect 245331 476307 245397 476308
rect 246438 476237 246498 479710
rect 247542 476237 247602 479710
rect 248278 476645 248338 479710
rect 248275 476644 248341 476645
rect 248275 476580 248276 476644
rect 248340 476580 248341 476644
rect 248275 476579 248341 476580
rect 248646 476237 248706 479710
rect 250118 476237 250178 479710
rect 250670 479710 250804 479770
rect 251288 479770 251348 480080
rect 252376 479770 252436 480080
rect 253464 479770 253524 480080
rect 251288 479710 251466 479770
rect 250670 476509 250730 479710
rect 250667 476508 250733 476509
rect 250667 476444 250668 476508
rect 250732 476444 250733 476508
rect 250667 476443 250733 476444
rect 251406 476373 251466 479710
rect 252326 479710 252436 479770
rect 253430 479710 253524 479770
rect 253600 479770 253660 480080
rect 254552 479770 254612 480080
rect 255912 479770 255972 480080
rect 253600 479710 253674 479770
rect 251403 476372 251469 476373
rect 251403 476308 251404 476372
rect 251468 476308 251469 476372
rect 251403 476307 251469 476308
rect 252326 476237 252386 479710
rect 253430 476237 253490 479710
rect 253614 476645 253674 479710
rect 254534 479710 254612 479770
rect 255822 479710 255972 479770
rect 256048 479770 256108 480080
rect 257000 479770 257060 480080
rect 258088 479770 258148 480080
rect 258496 479770 258556 480080
rect 256048 479710 256250 479770
rect 257000 479710 257170 479770
rect 254534 477053 254594 479710
rect 254531 477052 254597 477053
rect 254531 476988 254532 477052
rect 254596 476988 254597 477052
rect 254531 476987 254597 476988
rect 253611 476644 253677 476645
rect 253611 476580 253612 476644
rect 253676 476580 253677 476644
rect 253611 476579 253677 476580
rect 255822 476237 255882 479710
rect 256190 476917 256250 479710
rect 256187 476916 256253 476917
rect 256187 476852 256188 476916
rect 256252 476852 256253 476916
rect 256187 476851 256253 476852
rect 257110 476237 257170 479710
rect 257846 479710 258148 479770
rect 258398 479710 258556 479770
rect 259448 479770 259508 480080
rect 260672 479770 260732 480080
rect 261080 479770 261140 480080
rect 261760 479770 261820 480080
rect 262848 479770 262908 480080
rect 259448 479710 259562 479770
rect 257846 476645 257906 479710
rect 258398 476645 258458 479710
rect 257843 476644 257909 476645
rect 257843 476580 257844 476644
rect 257908 476580 257909 476644
rect 257843 476579 257909 476580
rect 258395 476644 258461 476645
rect 258395 476580 258396 476644
rect 258460 476580 258461 476644
rect 258395 476579 258461 476580
rect 259502 476237 259562 479710
rect 260606 479710 260732 479770
rect 260974 479710 261140 479770
rect 261710 479710 261820 479770
rect 262814 479710 262908 479770
rect 263528 479770 263588 480080
rect 263936 479770 263996 480080
rect 263528 479710 263610 479770
rect 260606 476373 260666 479710
rect 260974 476781 261034 479710
rect 260971 476780 261037 476781
rect 260971 476716 260972 476780
rect 261036 476716 261037 476780
rect 260971 476715 261037 476716
rect 260603 476372 260669 476373
rect 260603 476308 260604 476372
rect 260668 476308 260669 476372
rect 260603 476307 260669 476308
rect 261710 476237 261770 479710
rect 262814 476237 262874 479710
rect 263550 476645 263610 479710
rect 263918 479710 263996 479770
rect 265296 479770 265356 480080
rect 265976 479770 266036 480080
rect 265296 479710 265450 479770
rect 263547 476644 263613 476645
rect 263547 476580 263548 476644
rect 263612 476580 263613 476644
rect 263547 476579 263613 476580
rect 263918 476237 263978 479710
rect 265390 476237 265450 479710
rect 265942 479710 266036 479770
rect 266384 479770 266444 480080
rect 267608 479770 267668 480080
rect 266384 479710 266554 479770
rect 265942 477053 266002 479710
rect 265939 477052 266005 477053
rect 265939 476988 265940 477052
rect 266004 476988 266005 477052
rect 265939 476987 266005 476988
rect 266494 476373 266554 479710
rect 267598 479710 267668 479770
rect 268288 479770 268348 480080
rect 268696 479770 268756 480080
rect 269784 479770 269844 480080
rect 271008 479770 271068 480080
rect 268288 479710 268394 479770
rect 268696 479710 268762 479770
rect 269784 479710 269866 479770
rect 266491 476372 266557 476373
rect 266491 476308 266492 476372
rect 266556 476308 266557 476372
rect 266491 476307 266557 476308
rect 267598 476237 267658 479710
rect 268334 476509 268394 479710
rect 268331 476508 268397 476509
rect 268331 476444 268332 476508
rect 268396 476444 268397 476508
rect 268331 476443 268397 476444
rect 268702 476237 268762 479710
rect 269806 476237 269866 479710
rect 270910 479710 271068 479770
rect 271144 479770 271204 480080
rect 272232 479770 272292 480080
rect 273320 479770 273380 480080
rect 273592 479770 273652 480080
rect 274408 479770 274468 480080
rect 271144 479710 271338 479770
rect 270910 477053 270970 479710
rect 270907 477052 270973 477053
rect 270907 476988 270908 477052
rect 270972 476988 270973 477052
rect 270907 476987 270973 476988
rect 271278 476237 271338 479710
rect 272198 479710 272292 479770
rect 273302 479710 273380 479770
rect 273486 479710 273652 479770
rect 274406 479710 274468 479770
rect 275768 479770 275828 480080
rect 276040 479770 276100 480080
rect 276992 479770 277052 480080
rect 275768 479710 275938 479770
rect 276040 479710 276122 479770
rect 272198 476237 272258 479710
rect 273302 476373 273362 479710
rect 273486 476509 273546 479710
rect 273483 476508 273549 476509
rect 273483 476444 273484 476508
rect 273548 476444 273549 476508
rect 273483 476443 273549 476444
rect 273299 476372 273365 476373
rect 273299 476308 273300 476372
rect 273364 476308 273365 476372
rect 273299 476307 273365 476308
rect 274406 476237 274466 479710
rect 275878 476237 275938 479710
rect 276062 476645 276122 479710
rect 276982 479710 277052 479770
rect 278080 479770 278140 480080
rect 278488 479770 278548 480080
rect 278080 479710 278146 479770
rect 276059 476644 276125 476645
rect 276059 476580 276060 476644
rect 276124 476580 276125 476644
rect 276059 476579 276125 476580
rect 276982 476237 277042 479710
rect 278086 476237 278146 479710
rect 278454 479710 278548 479770
rect 279168 479770 279228 480080
rect 280936 479770 280996 480080
rect 283520 479770 283580 480080
rect 279168 479710 279250 479770
rect 278454 476917 278514 479710
rect 278451 476916 278517 476917
rect 278451 476852 278452 476916
rect 278516 476852 278517 476916
rect 278451 476851 278517 476852
rect 279190 476237 279250 479710
rect 280846 479710 280996 479770
rect 283422 479710 283580 479770
rect 285968 479770 286028 480080
rect 288280 479770 288340 480080
rect 291000 479770 291060 480080
rect 293448 479770 293508 480080
rect 285968 479710 286058 479770
rect 280846 476237 280906 479710
rect 283422 476237 283482 479710
rect 285998 476237 286058 479710
rect 288206 479710 288340 479770
rect 290966 479710 291060 479770
rect 293358 479710 293508 479770
rect 295896 479770 295956 480080
rect 298480 479770 298540 480080
rect 300928 479770 300988 480080
rect 303512 479770 303572 480080
rect 305960 479770 306020 480080
rect 308544 479770 308604 480080
rect 295896 479710 295994 479770
rect 298480 479710 298570 479770
rect 288206 476237 288266 479710
rect 290966 476237 291026 479710
rect 293358 476237 293418 479710
rect 295934 476237 295994 479710
rect 298510 476237 298570 479710
rect 300902 479710 300988 479770
rect 303478 479710 303572 479770
rect 305870 479710 306020 479770
rect 308446 479710 308604 479770
rect 310992 479770 311052 480080
rect 313440 479770 313500 480080
rect 315888 479770 315948 480080
rect 318472 479770 318532 480080
rect 310992 479710 311082 479770
rect 300902 476237 300962 479710
rect 303478 476781 303538 479710
rect 305870 477053 305930 479710
rect 308446 477053 308506 479710
rect 305867 477052 305933 477053
rect 305867 476988 305868 477052
rect 305932 476988 305933 477052
rect 305867 476987 305933 476988
rect 308443 477052 308509 477053
rect 308443 476988 308444 477052
rect 308508 476988 308509 477052
rect 308443 476987 308509 476988
rect 311022 476917 311082 479710
rect 313414 479710 313500 479770
rect 315806 479710 315948 479770
rect 318382 479710 318532 479770
rect 320920 479770 320980 480080
rect 323368 479770 323428 480080
rect 325952 479770 326012 480080
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 320920 479710 321018 479770
rect 311019 476916 311085 476917
rect 311019 476852 311020 476916
rect 311084 476852 311085 476916
rect 311019 476851 311085 476852
rect 303475 476780 303541 476781
rect 303475 476716 303476 476780
rect 303540 476716 303541 476780
rect 303475 476715 303541 476716
rect 313414 476509 313474 479710
rect 315806 476509 315866 479710
rect 313411 476508 313477 476509
rect 313411 476444 313412 476508
rect 313476 476444 313477 476508
rect 313411 476443 313477 476444
rect 315803 476508 315869 476509
rect 315803 476444 315804 476508
rect 315868 476444 315869 476508
rect 315803 476443 315869 476444
rect 318382 476373 318442 479710
rect 320958 476373 321018 479710
rect 323350 479710 323428 479770
rect 325926 479710 326012 479770
rect 323350 476917 323410 479710
rect 323347 476916 323413 476917
rect 323347 476852 323348 476916
rect 323412 476852 323413 476916
rect 323347 476851 323413 476852
rect 318379 476372 318445 476373
rect 318379 476308 318380 476372
rect 318444 476308 318445 476372
rect 318379 476307 318445 476308
rect 320955 476372 321021 476373
rect 320955 476308 320956 476372
rect 321020 476308 321021 476372
rect 320955 476307 321021 476308
rect 325926 476237 325986 479710
rect 235947 476236 236013 476237
rect 235947 476172 235948 476236
rect 236012 476172 236013 476236
rect 235947 476171 236013 476172
rect 238155 476236 238221 476237
rect 238155 476172 238156 476236
rect 238220 476172 238221 476236
rect 238155 476171 238221 476172
rect 239627 476236 239693 476237
rect 239627 476172 239628 476236
rect 239692 476172 239693 476236
rect 239627 476171 239693 476172
rect 240547 476236 240613 476237
rect 240547 476172 240548 476236
rect 240612 476172 240613 476236
rect 240547 476171 240613 476172
rect 241835 476236 241901 476237
rect 241835 476172 241836 476236
rect 241900 476172 241901 476236
rect 241835 476171 241901 476172
rect 246435 476236 246501 476237
rect 246435 476172 246436 476236
rect 246500 476172 246501 476236
rect 246435 476171 246501 476172
rect 247539 476236 247605 476237
rect 247539 476172 247540 476236
rect 247604 476172 247605 476236
rect 247539 476171 247605 476172
rect 248643 476236 248709 476237
rect 248643 476172 248644 476236
rect 248708 476172 248709 476236
rect 248643 476171 248709 476172
rect 250115 476236 250181 476237
rect 250115 476172 250116 476236
rect 250180 476172 250181 476236
rect 250115 476171 250181 476172
rect 252323 476236 252389 476237
rect 252323 476172 252324 476236
rect 252388 476172 252389 476236
rect 252323 476171 252389 476172
rect 253427 476236 253493 476237
rect 253427 476172 253428 476236
rect 253492 476172 253493 476236
rect 253427 476171 253493 476172
rect 255819 476236 255885 476237
rect 255819 476172 255820 476236
rect 255884 476172 255885 476236
rect 255819 476171 255885 476172
rect 257107 476236 257173 476237
rect 257107 476172 257108 476236
rect 257172 476172 257173 476236
rect 257107 476171 257173 476172
rect 259499 476236 259565 476237
rect 259499 476172 259500 476236
rect 259564 476172 259565 476236
rect 259499 476171 259565 476172
rect 261707 476236 261773 476237
rect 261707 476172 261708 476236
rect 261772 476172 261773 476236
rect 261707 476171 261773 476172
rect 262811 476236 262877 476237
rect 262811 476172 262812 476236
rect 262876 476172 262877 476236
rect 262811 476171 262877 476172
rect 263915 476236 263981 476237
rect 263915 476172 263916 476236
rect 263980 476172 263981 476236
rect 263915 476171 263981 476172
rect 265387 476236 265453 476237
rect 265387 476172 265388 476236
rect 265452 476172 265453 476236
rect 265387 476171 265453 476172
rect 267595 476236 267661 476237
rect 267595 476172 267596 476236
rect 267660 476172 267661 476236
rect 267595 476171 267661 476172
rect 268699 476236 268765 476237
rect 268699 476172 268700 476236
rect 268764 476172 268765 476236
rect 268699 476171 268765 476172
rect 269803 476236 269869 476237
rect 269803 476172 269804 476236
rect 269868 476172 269869 476236
rect 269803 476171 269869 476172
rect 271275 476236 271341 476237
rect 271275 476172 271276 476236
rect 271340 476172 271341 476236
rect 271275 476171 271341 476172
rect 272195 476236 272261 476237
rect 272195 476172 272196 476236
rect 272260 476172 272261 476236
rect 272195 476171 272261 476172
rect 274403 476236 274469 476237
rect 274403 476172 274404 476236
rect 274468 476172 274469 476236
rect 274403 476171 274469 476172
rect 275875 476236 275941 476237
rect 275875 476172 275876 476236
rect 275940 476172 275941 476236
rect 275875 476171 275941 476172
rect 276979 476236 277045 476237
rect 276979 476172 276980 476236
rect 277044 476172 277045 476236
rect 276979 476171 277045 476172
rect 278083 476236 278149 476237
rect 278083 476172 278084 476236
rect 278148 476172 278149 476236
rect 278083 476171 278149 476172
rect 279187 476236 279253 476237
rect 279187 476172 279188 476236
rect 279252 476172 279253 476236
rect 279187 476171 279253 476172
rect 280843 476236 280909 476237
rect 280843 476172 280844 476236
rect 280908 476172 280909 476236
rect 280843 476171 280909 476172
rect 283419 476236 283485 476237
rect 283419 476172 283420 476236
rect 283484 476172 283485 476236
rect 283419 476171 283485 476172
rect 285995 476236 286061 476237
rect 285995 476172 285996 476236
rect 286060 476172 286061 476236
rect 285995 476171 286061 476172
rect 288203 476236 288269 476237
rect 288203 476172 288204 476236
rect 288268 476172 288269 476236
rect 288203 476171 288269 476172
rect 290963 476236 291029 476237
rect 290963 476172 290964 476236
rect 291028 476172 291029 476236
rect 290963 476171 291029 476172
rect 293355 476236 293421 476237
rect 293355 476172 293356 476236
rect 293420 476172 293421 476236
rect 293355 476171 293421 476172
rect 295931 476236 295997 476237
rect 295931 476172 295932 476236
rect 295996 476172 295997 476236
rect 295931 476171 295997 476172
rect 298507 476236 298573 476237
rect 298507 476172 298508 476236
rect 298572 476172 298573 476236
rect 298507 476171 298573 476172
rect 300899 476236 300965 476237
rect 300899 476172 300900 476236
rect 300964 476172 300965 476236
rect 300899 476171 300965 476172
rect 325923 476236 325989 476237
rect 325923 476172 325924 476236
rect 325988 476172 325989 476236
rect 325923 476171 325989 476172
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 445423 362414 470898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 249568 439954 249888 439986
rect 249568 439718 249610 439954
rect 249846 439718 249888 439954
rect 249568 439634 249888 439718
rect 249568 439398 249610 439634
rect 249846 439398 249888 439634
rect 249568 439366 249888 439398
rect 280288 439954 280608 439986
rect 280288 439718 280330 439954
rect 280566 439718 280608 439954
rect 280288 439634 280608 439718
rect 280288 439398 280330 439634
rect 280566 439398 280608 439634
rect 280288 439366 280608 439398
rect 311008 439954 311328 439986
rect 311008 439718 311050 439954
rect 311286 439718 311328 439954
rect 311008 439634 311328 439718
rect 311008 439398 311050 439634
rect 311286 439398 311328 439634
rect 311008 439366 311328 439398
rect 341728 439954 342048 439986
rect 341728 439718 341770 439954
rect 342006 439718 342048 439954
rect 341728 439634 342048 439718
rect 341728 439398 341770 439634
rect 342006 439398 342048 439634
rect 341728 439366 342048 439398
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 234208 435454 234528 435486
rect 234208 435218 234250 435454
rect 234486 435218 234528 435454
rect 234208 435134 234528 435218
rect 234208 434898 234250 435134
rect 234486 434898 234528 435134
rect 234208 434866 234528 434898
rect 264928 435454 265248 435486
rect 264928 435218 264970 435454
rect 265206 435218 265248 435454
rect 264928 435134 265248 435218
rect 264928 434898 264970 435134
rect 265206 434898 265248 435134
rect 264928 434866 265248 434898
rect 295648 435454 295968 435486
rect 295648 435218 295690 435454
rect 295926 435218 295968 435454
rect 295648 435134 295968 435218
rect 295648 434898 295690 435134
rect 295926 434898 295968 435134
rect 295648 434866 295968 434898
rect 326368 435454 326688 435486
rect 326368 435218 326410 435454
rect 326646 435218 326688 435454
rect 326368 435134 326688 435218
rect 326368 434898 326410 435134
rect 326646 434898 326688 435134
rect 326368 434866 326688 434898
rect 357088 435454 357408 435486
rect 357088 435218 357130 435454
rect 357366 435218 357408 435454
rect 357088 435134 357408 435218
rect 357088 434898 357130 435134
rect 357366 434898 357408 435134
rect 357088 434866 357408 434898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 249568 403954 249888 403986
rect 249568 403718 249610 403954
rect 249846 403718 249888 403954
rect 249568 403634 249888 403718
rect 249568 403398 249610 403634
rect 249846 403398 249888 403634
rect 249568 403366 249888 403398
rect 280288 403954 280608 403986
rect 280288 403718 280330 403954
rect 280566 403718 280608 403954
rect 280288 403634 280608 403718
rect 280288 403398 280330 403634
rect 280566 403398 280608 403634
rect 280288 403366 280608 403398
rect 311008 403954 311328 403986
rect 311008 403718 311050 403954
rect 311286 403718 311328 403954
rect 311008 403634 311328 403718
rect 311008 403398 311050 403634
rect 311286 403398 311328 403634
rect 311008 403366 311328 403398
rect 341728 403954 342048 403986
rect 341728 403718 341770 403954
rect 342006 403718 342048 403954
rect 341728 403634 342048 403718
rect 341728 403398 341770 403634
rect 342006 403398 342048 403634
rect 341728 403366 342048 403398
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 234208 399454 234528 399486
rect 234208 399218 234250 399454
rect 234486 399218 234528 399454
rect 234208 399134 234528 399218
rect 234208 398898 234250 399134
rect 234486 398898 234528 399134
rect 234208 398866 234528 398898
rect 264928 399454 265248 399486
rect 264928 399218 264970 399454
rect 265206 399218 265248 399454
rect 264928 399134 265248 399218
rect 264928 398898 264970 399134
rect 265206 398898 265248 399134
rect 264928 398866 265248 398898
rect 295648 399454 295968 399486
rect 295648 399218 295690 399454
rect 295926 399218 295968 399454
rect 295648 399134 295968 399218
rect 295648 398898 295690 399134
rect 295926 398898 295968 399134
rect 295648 398866 295968 398898
rect 326368 399454 326688 399486
rect 326368 399218 326410 399454
rect 326646 399218 326688 399454
rect 326368 399134 326688 399218
rect 326368 398898 326410 399134
rect 326646 398898 326688 399134
rect 326368 398866 326688 398898
rect 357088 399454 357408 399486
rect 357088 399218 357130 399454
rect 357366 399218 357408 399454
rect 357088 399134 357408 399218
rect 357088 398898 357130 399134
rect 357366 398898 357408 399134
rect 357088 398866 357408 398898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 249568 367954 249888 367986
rect 249568 367718 249610 367954
rect 249846 367718 249888 367954
rect 249568 367634 249888 367718
rect 249568 367398 249610 367634
rect 249846 367398 249888 367634
rect 249568 367366 249888 367398
rect 280288 367954 280608 367986
rect 280288 367718 280330 367954
rect 280566 367718 280608 367954
rect 280288 367634 280608 367718
rect 280288 367398 280330 367634
rect 280566 367398 280608 367634
rect 280288 367366 280608 367398
rect 311008 367954 311328 367986
rect 311008 367718 311050 367954
rect 311286 367718 311328 367954
rect 311008 367634 311328 367718
rect 311008 367398 311050 367634
rect 311286 367398 311328 367634
rect 311008 367366 311328 367398
rect 341728 367954 342048 367986
rect 341728 367718 341770 367954
rect 342006 367718 342048 367954
rect 341728 367634 342048 367718
rect 341728 367398 341770 367634
rect 342006 367398 342048 367634
rect 341728 367366 342048 367398
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 234208 363454 234528 363486
rect 234208 363218 234250 363454
rect 234486 363218 234528 363454
rect 234208 363134 234528 363218
rect 234208 362898 234250 363134
rect 234486 362898 234528 363134
rect 234208 362866 234528 362898
rect 264928 363454 265248 363486
rect 264928 363218 264970 363454
rect 265206 363218 265248 363454
rect 264928 363134 265248 363218
rect 264928 362898 264970 363134
rect 265206 362898 265248 363134
rect 264928 362866 265248 362898
rect 295648 363454 295968 363486
rect 295648 363218 295690 363454
rect 295926 363218 295968 363454
rect 295648 363134 295968 363218
rect 295648 362898 295690 363134
rect 295926 362898 295968 363134
rect 295648 362866 295968 362898
rect 326368 363454 326688 363486
rect 326368 363218 326410 363454
rect 326646 363218 326688 363454
rect 326368 363134 326688 363218
rect 326368 362898 326410 363134
rect 326646 362898 326688 363134
rect 326368 362866 326688 362898
rect 357088 363454 357408 363486
rect 357088 363218 357130 363454
rect 357366 363218 357408 363454
rect 357088 363134 357408 363218
rect 357088 362898 357130 363134
rect 357366 362898 357408 363134
rect 357088 362866 357408 362898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 249568 331954 249888 331986
rect 249568 331718 249610 331954
rect 249846 331718 249888 331954
rect 249568 331634 249888 331718
rect 249568 331398 249610 331634
rect 249846 331398 249888 331634
rect 249568 331366 249888 331398
rect 280288 331954 280608 331986
rect 280288 331718 280330 331954
rect 280566 331718 280608 331954
rect 280288 331634 280608 331718
rect 280288 331398 280330 331634
rect 280566 331398 280608 331634
rect 280288 331366 280608 331398
rect 311008 331954 311328 331986
rect 311008 331718 311050 331954
rect 311286 331718 311328 331954
rect 311008 331634 311328 331718
rect 311008 331398 311050 331634
rect 311286 331398 311328 331634
rect 311008 331366 311328 331398
rect 341728 331954 342048 331986
rect 341728 331718 341770 331954
rect 342006 331718 342048 331954
rect 341728 331634 342048 331718
rect 341728 331398 341770 331634
rect 342006 331398 342048 331634
rect 341728 331366 342048 331398
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 234208 327454 234528 327486
rect 234208 327218 234250 327454
rect 234486 327218 234528 327454
rect 234208 327134 234528 327218
rect 234208 326898 234250 327134
rect 234486 326898 234528 327134
rect 234208 326866 234528 326898
rect 264928 327454 265248 327486
rect 264928 327218 264970 327454
rect 265206 327218 265248 327454
rect 264928 327134 265248 327218
rect 264928 326898 264970 327134
rect 265206 326898 265248 327134
rect 264928 326866 265248 326898
rect 295648 327454 295968 327486
rect 295648 327218 295690 327454
rect 295926 327218 295968 327454
rect 295648 327134 295968 327218
rect 295648 326898 295690 327134
rect 295926 326898 295968 327134
rect 295648 326866 295968 326898
rect 326368 327454 326688 327486
rect 326368 327218 326410 327454
rect 326646 327218 326688 327454
rect 326368 327134 326688 327218
rect 326368 326898 326410 327134
rect 326646 326898 326688 327134
rect 326368 326866 326688 326898
rect 357088 327454 357408 327486
rect 357088 327218 357130 327454
rect 357366 327218 357408 327454
rect 357088 327134 357408 327218
rect 357088 326898 357130 327134
rect 357366 326898 357408 327134
rect 357088 326866 357408 326898
rect 286179 308820 286245 308821
rect 286179 308756 286180 308820
rect 286244 308756 286245 308820
rect 286179 308755 286245 308756
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 245308 227414 263898
rect 231294 304954 231914 308400
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 245308 231914 268398
rect 240294 277954 240914 308400
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 100272 223954 100620 223986
rect 100272 223718 100328 223954
rect 100564 223718 100620 223954
rect 100272 223634 100620 223718
rect 100272 223398 100328 223634
rect 100564 223398 100620 223634
rect 100272 223366 100620 223398
rect 236000 223954 236348 223986
rect 236000 223718 236056 223954
rect 236292 223718 236348 223954
rect 236000 223634 236348 223718
rect 236000 223398 236056 223634
rect 236292 223398 236348 223634
rect 236000 223366 236348 223398
rect 100952 219454 101300 219486
rect 100952 219218 101008 219454
rect 101244 219218 101300 219454
rect 100952 219134 101300 219218
rect 100952 218898 101008 219134
rect 101244 218898 101300 219134
rect 100952 218866 101300 218898
rect 235320 219454 235668 219486
rect 235320 219218 235376 219454
rect 235612 219218 235668 219454
rect 235320 219134 235668 219218
rect 235320 218898 235376 219134
rect 235612 218898 235668 219134
rect 235320 218866 235668 218898
rect 100272 187954 100620 187986
rect 100272 187718 100328 187954
rect 100564 187718 100620 187954
rect 100272 187634 100620 187718
rect 100272 187398 100328 187634
rect 100564 187398 100620 187634
rect 100272 187366 100620 187398
rect 236000 187954 236348 187986
rect 236000 187718 236056 187954
rect 236292 187718 236348 187954
rect 236000 187634 236348 187718
rect 236000 187398 236056 187634
rect 236292 187398 236348 187634
rect 236000 187366 236348 187398
rect 100952 183454 101300 183486
rect 100952 183218 101008 183454
rect 101244 183218 101300 183454
rect 100952 183134 101300 183218
rect 100952 182898 101008 183134
rect 101244 182898 101300 183134
rect 100952 182866 101300 182898
rect 235320 183454 235668 183486
rect 235320 183218 235376 183454
rect 235612 183218 235668 183454
rect 235320 183134 235668 183218
rect 235320 182898 235376 183134
rect 235612 182898 235668 183134
rect 235320 182866 235668 182898
rect 116056 159490 116116 160106
rect 117144 159490 117204 160106
rect 118232 159490 118292 160106
rect 116056 159430 116226 159490
rect 116166 158677 116226 159430
rect 117086 159430 117204 159490
rect 118190 159430 118292 159490
rect 119592 159490 119652 160106
rect 120544 159490 120604 160106
rect 121768 159490 121828 160106
rect 123128 159490 123188 160106
rect 124216 159490 124276 160106
rect 125440 159490 125500 160106
rect 126528 159490 126588 160106
rect 127616 159490 127676 160106
rect 119592 159430 119722 159490
rect 120544 159430 120642 159490
rect 121768 159430 121930 159490
rect 123128 159430 123218 159490
rect 124216 159430 124322 159490
rect 117086 158677 117146 159430
rect 116163 158676 116229 158677
rect 116163 158612 116164 158676
rect 116228 158612 116229 158676
rect 116163 158611 116229 158612
rect 117083 158676 117149 158677
rect 117083 158612 117084 158676
rect 117148 158612 117149 158676
rect 117083 158611 117149 158612
rect 118190 158405 118250 159430
rect 119662 158677 119722 159430
rect 120582 158677 120642 159430
rect 121870 158677 121930 159430
rect 123158 158677 123218 159430
rect 119659 158676 119725 158677
rect 119659 158612 119660 158676
rect 119724 158612 119725 158676
rect 119659 158611 119725 158612
rect 120579 158676 120645 158677
rect 120579 158612 120580 158676
rect 120644 158612 120645 158676
rect 120579 158611 120645 158612
rect 121867 158676 121933 158677
rect 121867 158612 121868 158676
rect 121932 158612 121933 158676
rect 121867 158611 121933 158612
rect 123155 158676 123221 158677
rect 123155 158612 123156 158676
rect 123220 158612 123221 158676
rect 123155 158611 123221 158612
rect 118187 158404 118253 158405
rect 118187 158340 118188 158404
rect 118252 158340 118253 158404
rect 118187 158339 118253 158340
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 138454 101414 158000
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 142954 105914 158000
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 147454 110414 158000
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 151954 114914 158000
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 156454 119414 158000
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 120454 119414 155898
rect 118794 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 119414 120454
rect 118794 120134 119414 120218
rect 118794 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 119414 120134
rect 118794 84454 119414 119898
rect 118794 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 119414 84454
rect 118794 84134 119414 84218
rect 118794 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 119414 84134
rect 118794 48454 119414 83898
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 124954 123914 158000
rect 124262 157589 124322 159430
rect 125366 159430 125500 159490
rect 126470 159430 126588 159490
rect 127574 159430 127676 159490
rect 128296 159490 128356 160106
rect 128704 159490 128764 160106
rect 128296 159430 128370 159490
rect 124259 157588 124325 157589
rect 124259 157524 124260 157588
rect 124324 157524 124325 157588
rect 124259 157523 124325 157524
rect 125366 157453 125426 159430
rect 126470 158677 126530 159430
rect 127574 158677 127634 159430
rect 128310 158813 128370 159430
rect 128678 159430 128764 159490
rect 130064 159490 130124 160106
rect 130744 159490 130804 160106
rect 131288 159490 131348 160106
rect 132376 159490 132436 160106
rect 133464 159490 133524 160106
rect 130064 159430 130210 159490
rect 128307 158812 128373 158813
rect 128307 158748 128308 158812
rect 128372 158748 128373 158812
rect 128307 158747 128373 158748
rect 128678 158677 128738 159430
rect 130150 158677 130210 159430
rect 130702 159430 130804 159490
rect 131254 159430 131348 159490
rect 132358 159430 132436 159490
rect 133462 159430 133524 159490
rect 133600 159490 133660 160106
rect 134552 159490 134612 160106
rect 135912 159490 135972 160106
rect 136048 159490 136108 160106
rect 137000 159490 137060 160106
rect 138088 159490 138148 160106
rect 133600 159430 133706 159490
rect 134552 159430 134626 159490
rect 126467 158676 126533 158677
rect 126467 158612 126468 158676
rect 126532 158612 126533 158676
rect 126467 158611 126533 158612
rect 127571 158676 127637 158677
rect 127571 158612 127572 158676
rect 127636 158612 127637 158676
rect 127571 158611 127637 158612
rect 128675 158676 128741 158677
rect 128675 158612 128676 158676
rect 128740 158612 128741 158676
rect 128675 158611 128741 158612
rect 130147 158676 130213 158677
rect 130147 158612 130148 158676
rect 130212 158612 130213 158676
rect 130147 158611 130213 158612
rect 125363 157452 125429 157453
rect 125363 157388 125364 157452
rect 125428 157388 125429 157452
rect 125363 157387 125429 157388
rect 123294 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 123914 124954
rect 123294 124634 123914 124718
rect 123294 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 123914 124634
rect 123294 88954 123914 124398
rect 123294 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 123914 88954
rect 123294 88634 123914 88718
rect 123294 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 123914 88634
rect 123294 52954 123914 88398
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 129454 128414 158000
rect 130702 157725 130762 159430
rect 131254 158677 131314 159430
rect 132358 158677 132418 159430
rect 133462 158677 133522 159430
rect 131251 158676 131317 158677
rect 131251 158612 131252 158676
rect 131316 158612 131317 158676
rect 131251 158611 131317 158612
rect 132355 158676 132421 158677
rect 132355 158612 132356 158676
rect 132420 158612 132421 158676
rect 132355 158611 132421 158612
rect 133459 158676 133525 158677
rect 133459 158612 133460 158676
rect 133524 158612 133525 158676
rect 133459 158611 133525 158612
rect 133646 158133 133706 159430
rect 134566 158677 134626 159430
rect 135854 159430 135972 159490
rect 136038 159430 136108 159490
rect 136958 159430 137060 159490
rect 138062 159430 138148 159490
rect 138496 159490 138556 160106
rect 139448 159490 139508 160106
rect 140672 159490 140732 160106
rect 138496 159430 138674 159490
rect 139448 159430 139594 159490
rect 134563 158676 134629 158677
rect 134563 158612 134564 158676
rect 134628 158612 134629 158676
rect 134563 158611 134629 158612
rect 135854 158541 135914 159430
rect 135851 158540 135917 158541
rect 135851 158476 135852 158540
rect 135916 158476 135917 158540
rect 135851 158475 135917 158476
rect 133643 158132 133709 158133
rect 133643 158068 133644 158132
rect 133708 158068 133709 158132
rect 133643 158067 133709 158068
rect 130699 157724 130765 157725
rect 130699 157660 130700 157724
rect 130764 157660 130765 157724
rect 130699 157659 130765 157660
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 133954 132914 158000
rect 136038 157861 136098 159430
rect 136958 158541 137018 159430
rect 138062 158541 138122 159430
rect 136955 158540 137021 158541
rect 136955 158476 136956 158540
rect 137020 158476 137021 158540
rect 136955 158475 137021 158476
rect 138059 158540 138125 158541
rect 138059 158476 138060 158540
rect 138124 158476 138125 158540
rect 138059 158475 138125 158476
rect 136035 157860 136101 157861
rect 136035 157796 136036 157860
rect 136100 157796 136101 157860
rect 136035 157795 136101 157796
rect 132294 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 132914 133954
rect 132294 133634 132914 133718
rect 132294 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 132914 133634
rect 132294 97954 132914 133398
rect 132294 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 132914 97954
rect 132294 97634 132914 97718
rect 132294 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 132914 97634
rect 132294 61954 132914 97398
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 138454 137414 158000
rect 138614 157453 138674 159430
rect 139534 157861 139594 159430
rect 140638 159430 140732 159490
rect 141080 159490 141140 160106
rect 141760 159490 141820 160106
rect 142848 159490 142908 160106
rect 141080 159430 141250 159490
rect 140638 157997 140698 159430
rect 141190 158269 141250 159430
rect 141742 159430 141820 159490
rect 142846 159430 142908 159490
rect 143528 159490 143588 160106
rect 143936 159490 143996 160106
rect 145296 159490 145356 160106
rect 145976 159490 146036 160106
rect 146384 159490 146444 160106
rect 143528 159430 143642 159490
rect 143936 159430 144010 159490
rect 141742 158269 141802 159430
rect 141187 158268 141253 158269
rect 141187 158204 141188 158268
rect 141252 158204 141253 158268
rect 141187 158203 141253 158204
rect 141739 158268 141805 158269
rect 141739 158204 141740 158268
rect 141804 158204 141805 158268
rect 141739 158203 141805 158204
rect 140635 157996 140701 157997
rect 140635 157932 140636 157996
rect 140700 157932 140701 157996
rect 140635 157931 140701 157932
rect 139531 157860 139597 157861
rect 139531 157796 139532 157860
rect 139596 157796 139597 157860
rect 139531 157795 139597 157796
rect 138611 157452 138677 157453
rect 138611 157388 138612 157452
rect 138676 157388 138677 157452
rect 138611 157387 138677 157388
rect 136794 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 137414 138454
rect 136794 138134 137414 138218
rect 136794 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 137414 138134
rect 136794 102454 137414 137898
rect 136794 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 137414 102454
rect 136794 102134 137414 102218
rect 136794 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 137414 102134
rect 136794 66454 137414 101898
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 142954 141914 158000
rect 142846 157589 142906 159430
rect 142843 157588 142909 157589
rect 142843 157524 142844 157588
rect 142908 157524 142909 157588
rect 142843 157523 142909 157524
rect 143582 157453 143642 159430
rect 143950 158269 144010 159430
rect 145238 159430 145356 159490
rect 145974 159430 146036 159490
rect 146342 159430 146444 159490
rect 147608 159490 147668 160106
rect 148288 159490 148348 160106
rect 148696 159490 148756 160106
rect 149784 159490 149844 160106
rect 151008 159490 151068 160106
rect 147608 159430 147690 159490
rect 148288 159430 148426 159490
rect 148696 159430 148794 159490
rect 149784 159430 149898 159490
rect 143947 158268 144013 158269
rect 143947 158204 143948 158268
rect 144012 158204 144013 158268
rect 143947 158203 144013 158204
rect 145238 157861 145298 159430
rect 145974 158269 146034 159430
rect 146342 158269 146402 159430
rect 145971 158268 146037 158269
rect 145971 158204 145972 158268
rect 146036 158204 146037 158268
rect 145971 158203 146037 158204
rect 146339 158268 146405 158269
rect 146339 158204 146340 158268
rect 146404 158204 146405 158268
rect 146339 158203 146405 158204
rect 145235 157860 145301 157861
rect 145235 157796 145236 157860
rect 145300 157796 145301 157860
rect 145235 157795 145301 157796
rect 143579 157452 143645 157453
rect 143579 157388 143580 157452
rect 143644 157388 143645 157452
rect 143579 157387 143645 157388
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 106954 141914 142398
rect 141294 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 141914 106954
rect 141294 106634 141914 106718
rect 141294 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 141914 106634
rect 141294 70954 141914 106398
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 147454 146414 158000
rect 147630 157861 147690 159430
rect 147627 157860 147693 157861
rect 147627 157796 147628 157860
rect 147692 157796 147693 157860
rect 147627 157795 147693 157796
rect 148366 157453 148426 159430
rect 148734 158541 148794 159430
rect 148731 158540 148797 158541
rect 148731 158476 148732 158540
rect 148796 158476 148797 158540
rect 148731 158475 148797 158476
rect 149838 157453 149898 159430
rect 150942 159430 151068 159490
rect 151144 159490 151204 160106
rect 152232 159490 152292 160106
rect 151144 159430 151370 159490
rect 150942 158269 151002 159430
rect 150939 158268 151005 158269
rect 150939 158204 150940 158268
rect 151004 158204 151005 158268
rect 150939 158203 151005 158204
rect 148363 157452 148429 157453
rect 148363 157388 148364 157452
rect 148428 157388 148429 157452
rect 148363 157387 148429 157388
rect 149835 157452 149901 157453
rect 149835 157388 149836 157452
rect 149900 157388 149901 157452
rect 149835 157387 149901 157388
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 151954 150914 158000
rect 151310 157453 151370 159430
rect 152230 159430 152292 159490
rect 153320 159490 153380 160106
rect 153592 159490 153652 160106
rect 154408 159490 154468 160106
rect 155768 159490 155828 160106
rect 156040 159629 156100 160106
rect 156037 159628 156103 159629
rect 156037 159564 156038 159628
rect 156102 159564 156103 159628
rect 156037 159563 156103 159564
rect 153320 159430 153394 159490
rect 153592 159430 153762 159490
rect 154408 159430 154498 159490
rect 152230 157453 152290 159430
rect 153334 157453 153394 159430
rect 153702 158949 153762 159430
rect 153699 158948 153765 158949
rect 153699 158884 153700 158948
rect 153764 158884 153765 158948
rect 153699 158883 153765 158884
rect 154438 157453 154498 159430
rect 155726 159430 155828 159490
rect 156992 159490 157052 160106
rect 158080 159490 158140 160106
rect 158488 159901 158548 160106
rect 158485 159900 158551 159901
rect 158485 159836 158486 159900
rect 158550 159836 158551 159900
rect 158485 159835 158551 159836
rect 159168 159490 159228 160106
rect 160936 159490 160996 160106
rect 156992 159430 157074 159490
rect 158080 159430 158178 159490
rect 159168 159430 159282 159490
rect 151307 157452 151373 157453
rect 151307 157388 151308 157452
rect 151372 157388 151373 157452
rect 151307 157387 151373 157388
rect 152227 157452 152293 157453
rect 152227 157388 152228 157452
rect 152292 157388 152293 157452
rect 152227 157387 152293 157388
rect 153331 157452 153397 157453
rect 153331 157388 153332 157452
rect 153396 157388 153397 157452
rect 153331 157387 153397 157388
rect 154435 157452 154501 157453
rect 154435 157388 154436 157452
rect 154500 157388 154501 157452
rect 154435 157387 154501 157388
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 115954 150914 151398
rect 150294 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 150914 115954
rect 150294 115634 150914 115718
rect 150294 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 150914 115634
rect 150294 79954 150914 115398
rect 150294 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 150914 79954
rect 150294 79634 150914 79718
rect 150294 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 150914 79634
rect 150294 43954 150914 79398
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 156454 155414 158000
rect 155726 157453 155786 159430
rect 157014 157453 157074 159430
rect 158118 158677 158178 159430
rect 159222 158677 159282 159430
rect 160878 159430 160996 159490
rect 163520 159490 163580 160106
rect 165968 159901 166028 160106
rect 165965 159900 166031 159901
rect 165965 159836 165966 159900
rect 166030 159836 166031 159900
rect 165965 159835 166031 159836
rect 168280 159490 168340 160106
rect 171000 159490 171060 160106
rect 173448 159901 173508 160106
rect 173445 159900 173511 159901
rect 173445 159836 173446 159900
rect 173510 159836 173511 159900
rect 173445 159835 173511 159836
rect 163520 159430 163698 159490
rect 160878 158677 160938 159430
rect 163638 159085 163698 159430
rect 168238 159430 168340 159490
rect 170998 159430 171060 159490
rect 175896 159490 175956 160106
rect 178480 159490 178540 160106
rect 180928 159490 180988 160106
rect 183512 159490 183572 160106
rect 185960 159490 186020 160106
rect 175896 159430 176026 159490
rect 178480 159430 178602 159490
rect 180928 159430 180994 159490
rect 163635 159084 163701 159085
rect 163635 159020 163636 159084
rect 163700 159020 163701 159084
rect 163635 159019 163701 159020
rect 168238 158677 168298 159430
rect 158115 158676 158181 158677
rect 158115 158612 158116 158676
rect 158180 158612 158181 158676
rect 158115 158611 158181 158612
rect 159219 158676 159285 158677
rect 159219 158612 159220 158676
rect 159284 158612 159285 158676
rect 159219 158611 159285 158612
rect 160875 158676 160941 158677
rect 160875 158612 160876 158676
rect 160940 158612 160941 158676
rect 160875 158611 160941 158612
rect 168235 158676 168301 158677
rect 168235 158612 168236 158676
rect 168300 158612 168301 158676
rect 168235 158611 168301 158612
rect 170998 158133 171058 159430
rect 170995 158132 171061 158133
rect 170995 158068 170996 158132
rect 171060 158068 171061 158132
rect 170995 158067 171061 158068
rect 155723 157452 155789 157453
rect 155723 157388 155724 157452
rect 155788 157388 155789 157452
rect 155723 157387 155789 157388
rect 157011 157452 157077 157453
rect 157011 157388 157012 157452
rect 157076 157388 157077 157452
rect 157011 157387 157077 157388
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 120454 155414 155898
rect 154794 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 155414 120454
rect 154794 120134 155414 120218
rect 154794 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 155414 120134
rect 154794 84454 155414 119898
rect 154794 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 155414 84454
rect 154794 84134 155414 84218
rect 154794 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 155414 84134
rect 154794 48454 155414 83898
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 124954 159914 158000
rect 159294 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 159914 124954
rect 159294 124634 159914 124718
rect 159294 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 159914 124634
rect 159294 88954 159914 124398
rect 159294 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 159914 88954
rect 159294 88634 159914 88718
rect 159294 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 159914 88634
rect 159294 52954 159914 88398
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 129454 164414 158000
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 133954 168914 158000
rect 168294 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 168914 133954
rect 168294 133634 168914 133718
rect 168294 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 168914 133634
rect 168294 97954 168914 133398
rect 168294 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 168914 97954
rect 168294 97634 168914 97718
rect 168294 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 168914 97634
rect 168294 61954 168914 97398
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 138454 173414 158000
rect 175966 157453 176026 159430
rect 178542 158405 178602 159430
rect 180934 158405 180994 159430
rect 183510 159430 183572 159490
rect 185902 159430 186020 159490
rect 188544 159490 188604 160106
rect 190992 159490 191052 160106
rect 193440 159490 193500 160106
rect 195888 159490 195948 160106
rect 198472 159490 198532 160106
rect 188544 159430 188722 159490
rect 190992 159430 191114 159490
rect 193440 159430 193506 159490
rect 183510 158405 183570 159430
rect 178539 158404 178605 158405
rect 178539 158340 178540 158404
rect 178604 158340 178605 158404
rect 178539 158339 178605 158340
rect 180931 158404 180997 158405
rect 180931 158340 180932 158404
rect 180996 158340 180997 158404
rect 180931 158339 180997 158340
rect 183507 158404 183573 158405
rect 183507 158340 183508 158404
rect 183572 158340 183573 158404
rect 183507 158339 183573 158340
rect 185902 158269 185962 159430
rect 185899 158268 185965 158269
rect 185899 158204 185900 158268
rect 185964 158204 185965 158268
rect 185899 158203 185965 158204
rect 175963 157452 176029 157453
rect 175963 157388 175964 157452
rect 176028 157388 176029 157452
rect 175963 157387 176029 157388
rect 172794 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 173414 138454
rect 172794 138134 173414 138218
rect 172794 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 173414 138134
rect 172794 102454 173414 137898
rect 172794 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 173414 102454
rect 172794 102134 173414 102218
rect 172794 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 173414 102134
rect 172794 66454 173414 101898
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 142954 177914 158000
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 106954 177914 142398
rect 177294 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 177914 106954
rect 177294 106634 177914 106718
rect 177294 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 177914 106634
rect 177294 70954 177914 106398
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 147454 182414 158000
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 151954 186914 158000
rect 188662 157997 188722 159430
rect 191054 158405 191114 159430
rect 191051 158404 191117 158405
rect 191051 158340 191052 158404
rect 191116 158340 191117 158404
rect 191051 158339 191117 158340
rect 193446 158269 193506 159430
rect 195838 159430 195948 159490
rect 198414 159430 198532 159490
rect 200920 159490 200980 160106
rect 203368 159490 203428 160106
rect 205952 159629 206012 160106
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 205949 159628 206015 159629
rect 205949 159564 205950 159628
rect 206014 159564 206015 159628
rect 205949 159563 206015 159564
rect 200920 159430 201050 159490
rect 203368 159430 203442 159490
rect 195838 158541 195898 159430
rect 195835 158540 195901 158541
rect 195835 158476 195836 158540
rect 195900 158476 195901 158540
rect 195835 158475 195901 158476
rect 193443 158268 193509 158269
rect 193443 158204 193444 158268
rect 193508 158204 193509 158268
rect 193443 158203 193509 158204
rect 188659 157996 188725 157997
rect 188659 157932 188660 157996
rect 188724 157932 188725 157996
rect 188659 157931 188725 157932
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 115954 186914 151398
rect 186294 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 186914 115954
rect 186294 115634 186914 115718
rect 186294 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 186914 115634
rect 186294 79954 186914 115398
rect 186294 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 186914 79954
rect 186294 79634 186914 79718
rect 186294 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 186914 79634
rect 186294 43954 186914 79398
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 156454 191414 158000
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 120454 191414 155898
rect 190794 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 191414 120454
rect 190794 120134 191414 120218
rect 190794 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 191414 120134
rect 190794 84454 191414 119898
rect 190794 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 191414 84454
rect 190794 84134 191414 84218
rect 190794 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 191414 84134
rect 190794 48454 191414 83898
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 124954 195914 158000
rect 198414 157589 198474 159430
rect 198411 157588 198477 157589
rect 198411 157524 198412 157588
rect 198476 157524 198477 157588
rect 198411 157523 198477 157524
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 129454 200414 158000
rect 200990 157589 201050 159430
rect 203382 157589 203442 159430
rect 200987 157588 201053 157589
rect 200987 157524 200988 157588
rect 201052 157524 201053 157588
rect 200987 157523 201053 157524
rect 203379 157588 203445 157589
rect 203379 157524 203380 157588
rect 203444 157524 203445 157588
rect 203379 157523 203445 157524
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 133954 204914 158000
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 138454 209414 158000
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 142954 213914 158000
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 147454 218414 158000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 151954 222914 158000
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 156454 227414 158000
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 124954 231914 158000
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 129454 236414 158000
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 282454 245414 308400
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 286954 249914 308400
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 291454 254414 308400
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 295954 258914 308400
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 300454 263414 308400
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 304954 267914 308400
rect 270539 308276 270605 308277
rect 270539 308212 270540 308276
rect 270604 308212 270605 308276
rect 270539 308211 270605 308212
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 270542 152421 270602 308211
rect 271794 273454 272414 308400
rect 273299 308004 273365 308005
rect 273299 307940 273300 308004
rect 273364 307940 273365 308004
rect 273299 307939 273365 307940
rect 274587 308004 274653 308005
rect 274587 307940 274588 308004
rect 274652 307940 274653 308004
rect 274587 307939 274653 307940
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 270539 152420 270605 152421
rect 270539 152356 270540 152420
rect 270604 152356 270605 152420
rect 270539 152355 270605 152356
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 129454 272414 164898
rect 273302 138685 273362 307939
rect 273483 307868 273549 307869
rect 273483 307804 273484 307868
rect 273548 307804 273549 307868
rect 273483 307803 273549 307804
rect 273486 159357 273546 307803
rect 273483 159356 273549 159357
rect 273483 159292 273484 159356
rect 273548 159292 273549 159356
rect 273483 159291 273549 159292
rect 273299 138684 273365 138685
rect 273299 138620 273300 138684
rect 273364 138620 273365 138684
rect 273299 138619 273365 138620
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 274590 127669 274650 307939
rect 274771 307868 274837 307869
rect 274771 307804 274772 307868
rect 274836 307804 274837 307868
rect 274771 307803 274837 307804
rect 274774 146981 274834 307803
rect 276294 277954 276914 308400
rect 277347 307868 277413 307869
rect 277347 307804 277348 307868
rect 277412 307804 277413 307868
rect 277347 307803 277413 307804
rect 278819 307868 278885 307869
rect 278819 307804 278820 307868
rect 278884 307804 278885 307868
rect 278819 307803 278885 307804
rect 280291 307868 280357 307869
rect 280291 307804 280292 307868
rect 280356 307804 280357 307868
rect 280291 307803 280357 307804
rect 277350 302250 277410 307803
rect 278635 306236 278701 306237
rect 278635 306172 278636 306236
rect 278700 306172 278701 306236
rect 278635 306171 278701 306172
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 277166 302190 277410 302250
rect 277166 175949 277226 302190
rect 277163 175948 277229 175949
rect 277163 175884 277164 175948
rect 277228 175884 277229 175948
rect 277163 175883 277229 175884
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 274771 146980 274837 146981
rect 274771 146916 274772 146980
rect 274836 146916 274837 146980
rect 274771 146915 274837 146916
rect 276294 133954 276914 169398
rect 278638 158677 278698 306171
rect 278635 158676 278701 158677
rect 278635 158612 278636 158676
rect 278700 158612 278701 158676
rect 278635 158611 278701 158612
rect 278822 151061 278882 307803
rect 279923 247756 279989 247757
rect 279923 247692 279924 247756
rect 279988 247692 279989 247756
rect 279923 247691 279989 247692
rect 278819 151060 278885 151061
rect 278819 150996 278820 151060
rect 278884 150996 278885 151060
rect 278819 150995 278885 150996
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 274587 127668 274653 127669
rect 274587 127604 274588 127668
rect 274652 127604 274653 127668
rect 274587 127603 274653 127604
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 279926 9485 279986 247691
rect 279923 9484 279989 9485
rect 279923 9420 279924 9484
rect 279988 9420 279989 9484
rect 279923 9419 279989 9420
rect 280294 3365 280354 307803
rect 280794 282454 281414 308400
rect 284707 308276 284773 308277
rect 284707 308212 284708 308276
rect 284772 308212 284773 308276
rect 284707 308211 284773 308212
rect 283419 308004 283485 308005
rect 283419 307940 283420 308004
rect 283484 307940 283485 308004
rect 283419 307939 283485 307940
rect 283051 307868 283117 307869
rect 283051 307804 283052 307868
rect 283116 307804 283117 307868
rect 283051 307803 283117 307804
rect 283054 302250 283114 307803
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 282870 302190 283114 302250
rect 282315 248028 282381 248029
rect 282315 247964 282316 248028
rect 282380 247964 282381 248028
rect 282315 247963 282381 247964
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280475 244900 280541 244901
rect 280475 244836 280476 244900
rect 280540 244836 280541 244900
rect 280475 244835 280541 244836
rect 280478 3909 280538 244835
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280475 3908 280541 3909
rect 280475 3844 280476 3908
rect 280540 3844 280541 3908
rect 280475 3843 280541 3844
rect 280291 3364 280357 3365
rect 280291 3300 280292 3364
rect 280356 3300 280357 3364
rect 280291 3299 280357 3300
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 -6106 281414 29898
rect 282318 9621 282378 247963
rect 282499 245036 282565 245037
rect 282499 244972 282500 245036
rect 282564 244972 282565 245036
rect 282499 244971 282565 244972
rect 282315 9620 282381 9621
rect 282315 9556 282316 9620
rect 282380 9556 282381 9620
rect 282315 9555 282381 9556
rect 282502 4045 282562 244971
rect 282683 244764 282749 244765
rect 282683 244700 282684 244764
rect 282748 244700 282749 244764
rect 282683 244699 282749 244700
rect 282499 4044 282565 4045
rect 282499 3980 282500 4044
rect 282564 3980 282565 4044
rect 282499 3979 282565 3980
rect 282686 3229 282746 244699
rect 282870 157350 282930 302190
rect 283422 158949 283482 307939
rect 283971 247620 284037 247621
rect 283971 247556 283972 247620
rect 284036 247556 284037 247620
rect 283971 247555 284037 247556
rect 283419 158948 283485 158949
rect 283419 158884 283420 158948
rect 283484 158884 283485 158948
rect 283419 158883 283485 158884
rect 282870 157290 283114 157350
rect 283054 147690 283114 157290
rect 282870 147630 283114 147690
rect 282870 125493 282930 147630
rect 282867 125492 282933 125493
rect 282867 125428 282868 125492
rect 282932 125428 282933 125492
rect 282867 125427 282933 125428
rect 283974 9213 284034 247555
rect 284155 247076 284221 247077
rect 284155 247012 284156 247076
rect 284220 247012 284221 247076
rect 284155 247011 284221 247012
rect 283971 9212 284037 9213
rect 283971 9148 283972 9212
rect 284036 9148 284037 9212
rect 283971 9147 284037 9148
rect 284158 8941 284218 247011
rect 284710 158813 284770 308211
rect 285294 286954 285914 308400
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285075 247892 285141 247893
rect 285075 247828 285076 247892
rect 285140 247828 285141 247892
rect 285075 247827 285141 247828
rect 284891 247076 284957 247077
rect 284891 247012 284892 247076
rect 284956 247012 284957 247076
rect 284891 247011 284957 247012
rect 284707 158812 284773 158813
rect 284707 158748 284708 158812
rect 284772 158748 284773 158812
rect 284707 158747 284773 158748
rect 284894 9077 284954 247011
rect 284891 9076 284957 9077
rect 284891 9012 284892 9076
rect 284956 9012 284957 9076
rect 284891 9011 284957 9012
rect 284155 8940 284221 8941
rect 284155 8876 284156 8940
rect 284220 8876 284221 8940
rect 284155 8875 284221 8876
rect 285078 3365 285138 247827
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 286182 159085 286242 308755
rect 292435 308684 292501 308685
rect 292435 308620 292436 308684
rect 292500 308620 292501 308684
rect 292435 308619 292501 308620
rect 297955 308684 298021 308685
rect 297955 308620 297956 308684
rect 298020 308620 298021 308684
rect 297955 308619 298021 308620
rect 287835 307868 287901 307869
rect 287835 307804 287836 307868
rect 287900 307804 287901 307868
rect 287835 307803 287901 307804
rect 286915 248164 286981 248165
rect 286915 248100 286916 248164
rect 286980 248100 286981 248164
rect 286915 248099 286981 248100
rect 286363 247076 286429 247077
rect 286363 247012 286364 247076
rect 286428 247012 286429 247076
rect 286363 247011 286429 247012
rect 286179 159084 286245 159085
rect 286179 159020 286180 159084
rect 286244 159020 286245 159084
rect 286179 159019 286245 159020
rect 286366 158813 286426 247011
rect 286731 245172 286797 245173
rect 286731 245108 286732 245172
rect 286796 245108 286797 245172
rect 286731 245107 286797 245108
rect 286363 158812 286429 158813
rect 286363 158748 286364 158812
rect 286428 158748 286429 158812
rect 286363 158747 286429 158748
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285075 3364 285141 3365
rect 285075 3300 285076 3364
rect 285140 3300 285141 3364
rect 285075 3299 285141 3300
rect 282683 3228 282749 3229
rect 282683 3164 282684 3228
rect 282748 3164 282749 3228
rect 282683 3163 282749 3164
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 -7066 285914 34398
rect 286734 6357 286794 245107
rect 286731 6356 286797 6357
rect 286731 6292 286732 6356
rect 286796 6292 286797 6356
rect 286731 6291 286797 6292
rect 286918 3637 286978 248099
rect 287651 247076 287717 247077
rect 287651 247012 287652 247076
rect 287716 247012 287717 247076
rect 287651 247011 287717 247012
rect 287654 158813 287714 247011
rect 287651 158812 287717 158813
rect 287651 158748 287652 158812
rect 287716 158748 287717 158812
rect 287651 158747 287717 158748
rect 287838 155277 287898 307803
rect 289794 291454 290414 308400
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 288203 248300 288269 248301
rect 288203 248236 288204 248300
rect 288268 248236 288269 248300
rect 288203 248235 288269 248236
rect 288019 244356 288085 244357
rect 288019 244292 288020 244356
rect 288084 244292 288085 244356
rect 288019 244291 288085 244292
rect 287835 155276 287901 155277
rect 287835 155212 287836 155276
rect 287900 155212 287901 155276
rect 287835 155211 287901 155212
rect 288022 6221 288082 244291
rect 288019 6220 288085 6221
rect 288019 6156 288020 6220
rect 288084 6156 288085 6220
rect 288019 6155 288085 6156
rect 286915 3636 286981 3637
rect 286915 3572 286916 3636
rect 286980 3572 286981 3636
rect 286915 3571 286981 3572
rect 288206 3501 288266 248235
rect 288755 247076 288821 247077
rect 288755 247012 288756 247076
rect 288820 247012 288821 247076
rect 288755 247011 288821 247012
rect 288758 158813 288818 247011
rect 289307 245580 289373 245581
rect 289307 245516 289308 245580
rect 289372 245516 289373 245580
rect 289307 245515 289373 245516
rect 289123 245444 289189 245445
rect 289123 245380 289124 245444
rect 289188 245380 289189 245444
rect 289123 245379 289189 245380
rect 288755 158812 288821 158813
rect 288755 158748 288756 158812
rect 288820 158748 288821 158812
rect 288755 158747 288821 158748
rect 289126 6629 289186 245379
rect 289310 6765 289370 245515
rect 289491 244628 289557 244629
rect 289491 244564 289492 244628
rect 289556 244564 289557 244628
rect 289491 244563 289557 244564
rect 289307 6764 289373 6765
rect 289307 6700 289308 6764
rect 289372 6700 289373 6764
rect 289307 6699 289373 6700
rect 289123 6628 289189 6629
rect 289123 6564 289124 6628
rect 289188 6564 289189 6628
rect 289123 6563 289189 6564
rect 289494 6493 289554 244563
rect 289794 219454 290414 254898
rect 292251 247484 292317 247485
rect 292251 247420 292252 247484
rect 292316 247420 292317 247484
rect 292251 247419 292317 247420
rect 290779 244492 290845 244493
rect 290779 244428 290780 244492
rect 290844 244428 290845 244492
rect 290779 244427 290845 244428
rect 290595 244356 290661 244357
rect 290595 244292 290596 244356
rect 290660 244292 290661 244356
rect 290595 244291 290661 244292
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 290598 158813 290658 244291
rect 290782 158813 290842 244427
rect 291699 244356 291765 244357
rect 291699 244292 291700 244356
rect 291764 244292 291765 244356
rect 291699 244291 291765 244292
rect 291883 244356 291949 244357
rect 291883 244292 291884 244356
rect 291948 244292 291949 244356
rect 291883 244291 291949 244292
rect 290595 158812 290661 158813
rect 290595 158748 290596 158812
rect 290660 158748 290661 158812
rect 290595 158747 290661 158748
rect 290779 158812 290845 158813
rect 290779 158748 290780 158812
rect 290844 158748 290845 158812
rect 290779 158747 290845 158748
rect 291702 157453 291762 244291
rect 291886 158813 291946 244291
rect 291883 158812 291949 158813
rect 291883 158748 291884 158812
rect 291948 158748 291949 158812
rect 291883 158747 291949 158748
rect 291699 157452 291765 157453
rect 291699 157388 291700 157452
rect 291764 157388 291765 157452
rect 291699 157387 291765 157388
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289491 6492 289557 6493
rect 289491 6428 289492 6492
rect 289556 6428 289557 6492
rect 289491 6427 289557 6428
rect 288203 3500 288269 3501
rect 288203 3436 288204 3500
rect 288268 3436 288269 3500
rect 288203 3435 288269 3436
rect 289794 3454 290414 38898
rect 292254 9349 292314 247419
rect 292251 9348 292317 9349
rect 292251 9284 292252 9348
rect 292316 9284 292317 9348
rect 292251 9283 292317 9284
rect 292438 8805 292498 308619
rect 293723 307868 293789 307869
rect 293723 307804 293724 307868
rect 293788 307804 293789 307868
rect 293723 307803 293789 307804
rect 293171 247076 293237 247077
rect 293171 247012 293172 247076
rect 293236 247012 293237 247076
rect 293171 247011 293237 247012
rect 293174 149157 293234 247011
rect 293539 245308 293605 245309
rect 293539 245244 293540 245308
rect 293604 245244 293605 245308
rect 293539 245243 293605 245244
rect 293355 244764 293421 244765
rect 293355 244700 293356 244764
rect 293420 244700 293421 244764
rect 293355 244699 293421 244700
rect 293358 158813 293418 244699
rect 293542 167109 293602 245243
rect 293539 167108 293605 167109
rect 293539 167044 293540 167108
rect 293604 167044 293605 167108
rect 293539 167043 293605 167044
rect 293355 158812 293421 158813
rect 293355 158748 293356 158812
rect 293420 158748 293421 158812
rect 293355 158747 293421 158748
rect 293171 149156 293237 149157
rect 293171 149092 293172 149156
rect 293236 149092 293237 149156
rect 293171 149091 293237 149092
rect 293726 148341 293786 307803
rect 294294 295954 294914 308400
rect 297771 308140 297837 308141
rect 297771 308076 297772 308140
rect 297836 308076 297837 308140
rect 297771 308075 297837 308076
rect 296299 307868 296365 307869
rect 296299 307804 296300 307868
rect 296364 307804 296365 307868
rect 296299 307803 296365 307804
rect 296483 307868 296549 307869
rect 296483 307804 296484 307868
rect 296548 307804 296549 307868
rect 296483 307803 296549 307804
rect 297587 307868 297653 307869
rect 297587 307804 297588 307868
rect 297652 307804 297653 307868
rect 297587 307803 297653 307804
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 295011 247076 295077 247077
rect 295011 247012 295012 247076
rect 295076 247012 295077 247076
rect 295011 247011 295077 247012
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 295014 158813 295074 247011
rect 296115 245444 296181 245445
rect 296115 245380 296116 245444
rect 296180 245380 296181 245444
rect 296115 245379 296181 245380
rect 295195 244900 295261 244901
rect 295195 244836 295196 244900
rect 295260 244836 295261 244900
rect 295195 244835 295261 244836
rect 295198 195261 295258 244835
rect 295931 244764 295997 244765
rect 295931 244700 295932 244764
rect 295996 244700 295997 244764
rect 295931 244699 295997 244700
rect 295195 195260 295261 195261
rect 295195 195196 295196 195260
rect 295260 195196 295261 195260
rect 295195 195195 295261 195196
rect 295934 158813 295994 244699
rect 295011 158812 295077 158813
rect 295011 158748 295012 158812
rect 295076 158748 295077 158812
rect 295011 158747 295077 158748
rect 295931 158812 295997 158813
rect 295931 158748 295932 158812
rect 295996 158748 295997 158812
rect 295931 158747 295997 158748
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 293723 148340 293789 148341
rect 293723 148276 293724 148340
rect 293788 148276 293789 148340
rect 293723 148275 293789 148276
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 292435 8804 292501 8805
rect 292435 8740 292436 8804
rect 292500 8740 292501 8804
rect 292435 8739 292501 8740
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 296118 3773 296178 245379
rect 296302 7581 296362 307803
rect 296299 7580 296365 7581
rect 296299 7516 296300 7580
rect 296364 7516 296365 7580
rect 296299 7515 296365 7516
rect 296486 4997 296546 307803
rect 297590 6085 297650 307803
rect 297774 6901 297834 308075
rect 297771 6900 297837 6901
rect 297771 6836 297772 6900
rect 297836 6836 297837 6900
rect 297771 6835 297837 6836
rect 297587 6084 297653 6085
rect 297587 6020 297588 6084
rect 297652 6020 297653 6084
rect 297587 6019 297653 6020
rect 296483 4996 296549 4997
rect 296483 4932 296484 4996
rect 296548 4932 296549 4996
rect 296483 4931 296549 4932
rect 297958 4861 298018 308619
rect 298323 308140 298389 308141
rect 298323 308076 298324 308140
rect 298388 308076 298389 308140
rect 298323 308075 298389 308076
rect 298139 245580 298205 245581
rect 298139 245516 298140 245580
rect 298204 245516 298205 245580
rect 298139 245515 298205 245516
rect 298142 152421 298202 245515
rect 298326 159357 298386 308075
rect 298507 307868 298573 307869
rect 298507 307804 298508 307868
rect 298572 307804 298573 307868
rect 298507 307803 298573 307804
rect 298323 159356 298389 159357
rect 298323 159292 298324 159356
rect 298388 159292 298389 159356
rect 298323 159291 298389 159292
rect 298139 152420 298205 152421
rect 298139 152356 298140 152420
rect 298204 152356 298205 152420
rect 298139 152355 298205 152356
rect 298510 82109 298570 307803
rect 298794 300454 299414 308400
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 245308 299414 263898
rect 303294 304954 303914 308400
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 245308 303914 268398
rect 316794 282454 317414 308400
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 245308 317414 245898
rect 321294 286954 321914 308400
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 245308 321914 250398
rect 325794 291454 326414 308400
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 245308 326414 254898
rect 330294 295954 330914 308400
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 245308 330914 259398
rect 334794 300454 335414 308400
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 245308 335414 263898
rect 339294 304954 339914 308400
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 245308 339914 268398
rect 352794 282454 353414 308400
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 245308 353414 245898
rect 357294 286954 357914 308400
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 245308 357914 250398
rect 361794 291454 362414 308400
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 245308 362414 254898
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 245308 366914 259398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 245308 371414 263898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 245308 375914 268398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 245308 380414 272898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 245308 384914 277398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 245308 389414 245898
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 245308 393914 250398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 245308 398414 254898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 245308 402914 259398
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 245308 407414 263898
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 245308 411914 268398
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 245308 416414 272898
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 245308 420914 277398
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 245308 425414 245898
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 245308 429914 250398
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 439451 444412 439517 444413
rect 439451 444348 439452 444412
rect 439516 444348 439517 444412
rect 439451 444347 439517 444348
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 437427 297396 437493 297397
rect 437427 297332 437428 297396
rect 437492 297332 437493 297396
rect 437427 297331 437493 297332
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 245308 434414 254898
rect 299059 245172 299125 245173
rect 299059 245108 299060 245172
rect 299124 245108 299125 245172
rect 299059 245107 299125 245108
rect 299062 196077 299122 245107
rect 300272 223954 300620 223986
rect 300272 223718 300328 223954
rect 300564 223718 300620 223954
rect 300272 223634 300620 223718
rect 300272 223398 300328 223634
rect 300564 223398 300620 223634
rect 300272 223366 300620 223398
rect 436000 223954 436348 223986
rect 436000 223718 436056 223954
rect 436292 223718 436348 223954
rect 436000 223634 436348 223718
rect 436000 223398 436056 223634
rect 436292 223398 436348 223634
rect 436000 223366 436348 223398
rect 300952 219454 301300 219486
rect 300952 219218 301008 219454
rect 301244 219218 301300 219454
rect 300952 219134 301300 219218
rect 300952 218898 301008 219134
rect 301244 218898 301300 219134
rect 300952 218866 301300 218898
rect 435320 219454 435668 219486
rect 435320 219218 435376 219454
rect 435612 219218 435668 219454
rect 435320 219134 435668 219218
rect 435320 218898 435376 219134
rect 435612 218898 435668 219134
rect 435320 218866 435668 218898
rect 299059 196076 299125 196077
rect 299059 196012 299060 196076
rect 299124 196012 299125 196076
rect 299059 196011 299125 196012
rect 300272 187954 300620 187986
rect 300272 187718 300328 187954
rect 300564 187718 300620 187954
rect 300272 187634 300620 187718
rect 300272 187398 300328 187634
rect 300564 187398 300620 187634
rect 300272 187366 300620 187398
rect 436000 187954 436348 187986
rect 436000 187718 436056 187954
rect 436292 187718 436348 187954
rect 436000 187634 436348 187718
rect 436000 187398 436056 187634
rect 436292 187398 436348 187634
rect 436000 187366 436348 187398
rect 300952 183454 301300 183486
rect 300952 183218 301008 183454
rect 301244 183218 301300 183454
rect 300952 183134 301300 183218
rect 300952 182898 301008 183134
rect 301244 182898 301300 183134
rect 300952 182866 301300 182898
rect 435320 183454 435668 183486
rect 435320 183218 435376 183454
rect 435612 183218 435668 183454
rect 435320 183134 435668 183218
rect 435320 182898 435376 183134
rect 435612 182898 435668 183134
rect 435320 182866 435668 182898
rect 316056 159490 316116 160106
rect 317144 159490 317204 160106
rect 318232 159490 318292 160106
rect 319592 159490 319652 160106
rect 315806 159430 316116 159490
rect 317094 159430 317204 159490
rect 318198 159430 318292 159490
rect 319486 159430 319652 159490
rect 320544 159490 320604 160106
rect 321768 159490 321828 160106
rect 320544 159430 320650 159490
rect 315806 158677 315866 159430
rect 317094 158677 317154 159430
rect 318198 158677 318258 159430
rect 319486 158677 319546 159430
rect 320590 158677 320650 159430
rect 321694 159430 321828 159490
rect 323128 159490 323188 160106
rect 324216 159490 324276 160106
rect 325440 159490 325500 160106
rect 326528 159490 326588 160106
rect 327616 159490 327676 160106
rect 323128 159430 323226 159490
rect 324216 159430 324330 159490
rect 321694 158677 321754 159430
rect 323166 158677 323226 159430
rect 315803 158676 315869 158677
rect 315803 158612 315804 158676
rect 315868 158612 315869 158676
rect 315803 158611 315869 158612
rect 317091 158676 317157 158677
rect 317091 158612 317092 158676
rect 317156 158612 317157 158676
rect 317091 158611 317157 158612
rect 318195 158676 318261 158677
rect 318195 158612 318196 158676
rect 318260 158612 318261 158676
rect 318195 158611 318261 158612
rect 319483 158676 319549 158677
rect 319483 158612 319484 158676
rect 319548 158612 319549 158676
rect 319483 158611 319549 158612
rect 320587 158676 320653 158677
rect 320587 158612 320588 158676
rect 320652 158612 320653 158676
rect 320587 158611 320653 158612
rect 321691 158676 321757 158677
rect 321691 158612 321692 158676
rect 321756 158612 321757 158676
rect 321691 158611 321757 158612
rect 323163 158676 323229 158677
rect 323163 158612 323164 158676
rect 323228 158612 323229 158676
rect 323163 158611 323229 158612
rect 298794 156454 299414 158000
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298507 82108 298573 82109
rect 298507 82044 298508 82108
rect 298572 82044 298573 82108
rect 298507 82043 298573 82044
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 297955 4860 298021 4861
rect 297955 4796 297956 4860
rect 298020 4796 298021 4860
rect 297955 4795 298021 4796
rect 296115 3772 296181 3773
rect 296115 3708 296116 3772
rect 296180 3708 296181 3772
rect 296115 3707 296181 3708
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 124954 303914 158000
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 129454 308414 158000
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 133954 312914 158000
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 138454 317414 158000
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 142954 321914 158000
rect 324270 157861 324330 159430
rect 325374 159430 325500 159490
rect 326478 159430 326588 159490
rect 327582 159430 327676 159490
rect 328296 159490 328356 160106
rect 328704 159490 328764 160106
rect 330064 159490 330124 160106
rect 330744 159490 330804 160106
rect 331288 159490 331348 160106
rect 332376 159490 332436 160106
rect 328296 159430 328378 159490
rect 324267 157860 324333 157861
rect 324267 157796 324268 157860
rect 324332 157796 324333 157860
rect 324267 157795 324333 157796
rect 325374 157453 325434 159430
rect 326478 158677 326538 159430
rect 326475 158676 326541 158677
rect 326475 158612 326476 158676
rect 326540 158612 326541 158676
rect 326475 158611 326541 158612
rect 325371 157452 325437 157453
rect 325371 157388 325372 157452
rect 325436 157388 325437 157452
rect 325371 157387 325437 157388
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 147454 326414 158000
rect 327582 157997 327642 159430
rect 328318 158677 328378 159430
rect 328686 159430 328764 159490
rect 329974 159430 330124 159490
rect 330710 159430 330804 159490
rect 331262 159430 331348 159490
rect 332366 159430 332436 159490
rect 333464 159490 333524 160106
rect 333600 159490 333660 160106
rect 334552 159490 334612 160106
rect 335912 159490 335972 160106
rect 336048 159901 336108 160106
rect 336045 159900 336111 159901
rect 336045 159836 336046 159900
rect 336110 159836 336111 159900
rect 336045 159835 336111 159836
rect 337000 159490 337060 160106
rect 338088 159490 338148 160106
rect 338496 159901 338556 160106
rect 338493 159900 338559 159901
rect 338493 159836 338494 159900
rect 338558 159836 338559 159900
rect 338493 159835 338559 159836
rect 339448 159490 339508 160106
rect 340672 159490 340732 160106
rect 341080 159490 341140 160106
rect 341760 159490 341820 160106
rect 333464 159430 333530 159490
rect 333600 159430 333714 159490
rect 334552 159430 334634 159490
rect 328315 158676 328381 158677
rect 328315 158612 328316 158676
rect 328380 158612 328381 158676
rect 328315 158611 328381 158612
rect 328686 158133 328746 159430
rect 329974 158677 330034 159430
rect 330710 158677 330770 159430
rect 329971 158676 330037 158677
rect 329971 158612 329972 158676
rect 330036 158612 330037 158676
rect 329971 158611 330037 158612
rect 330707 158676 330773 158677
rect 330707 158612 330708 158676
rect 330772 158612 330773 158676
rect 330707 158611 330773 158612
rect 331262 158269 331322 159430
rect 332366 158405 332426 159430
rect 333470 158677 333530 159430
rect 333467 158676 333533 158677
rect 333467 158612 333468 158676
rect 333532 158612 333533 158676
rect 333467 158611 333533 158612
rect 333654 158405 333714 159430
rect 334574 158677 334634 159430
rect 335862 159430 335972 159490
rect 336966 159430 337060 159490
rect 338070 159430 338148 159490
rect 339358 159430 339508 159490
rect 340646 159430 340732 159490
rect 341014 159430 341140 159490
rect 341750 159430 341820 159490
rect 342848 159490 342908 160106
rect 343528 159490 343588 160106
rect 343936 159490 343996 160106
rect 345296 159490 345356 160106
rect 342848 159430 342914 159490
rect 343528 159430 343650 159490
rect 343936 159430 344018 159490
rect 335862 158677 335922 159430
rect 334571 158676 334637 158677
rect 334571 158612 334572 158676
rect 334636 158612 334637 158676
rect 334571 158611 334637 158612
rect 335859 158676 335925 158677
rect 335859 158612 335860 158676
rect 335924 158612 335925 158676
rect 335859 158611 335925 158612
rect 336966 158405 337026 159430
rect 338070 158677 338130 159430
rect 338067 158676 338133 158677
rect 338067 158612 338068 158676
rect 338132 158612 338133 158676
rect 338067 158611 338133 158612
rect 332363 158404 332429 158405
rect 332363 158340 332364 158404
rect 332428 158340 332429 158404
rect 332363 158339 332429 158340
rect 333651 158404 333717 158405
rect 333651 158340 333652 158404
rect 333716 158340 333717 158404
rect 333651 158339 333717 158340
rect 336963 158404 337029 158405
rect 336963 158340 336964 158404
rect 337028 158340 337029 158404
rect 336963 158339 337029 158340
rect 339358 158269 339418 159430
rect 331259 158268 331325 158269
rect 331259 158204 331260 158268
rect 331324 158204 331325 158268
rect 331259 158203 331325 158204
rect 339355 158268 339421 158269
rect 339355 158204 339356 158268
rect 339420 158204 339421 158268
rect 339355 158203 339421 158204
rect 328683 158132 328749 158133
rect 328683 158068 328684 158132
rect 328748 158068 328749 158132
rect 328683 158067 328749 158068
rect 327579 157996 327645 157997
rect 327579 157932 327580 157996
rect 327644 157932 327645 157996
rect 327579 157931 327645 157932
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 151954 330914 158000
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 156454 335414 158000
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 124954 339914 158000
rect 340646 157997 340706 159430
rect 341014 158677 341074 159430
rect 341011 158676 341077 158677
rect 341011 158612 341012 158676
rect 341076 158612 341077 158676
rect 341011 158611 341077 158612
rect 340643 157996 340709 157997
rect 340643 157932 340644 157996
rect 340708 157932 340709 157996
rect 340643 157931 340709 157932
rect 341750 157861 341810 159430
rect 342854 157997 342914 159430
rect 343590 158677 343650 159430
rect 343958 158677 344018 159430
rect 345246 159430 345356 159490
rect 345976 159490 346036 160106
rect 346384 159490 346444 160106
rect 345976 159430 346042 159490
rect 343587 158676 343653 158677
rect 343587 158612 343588 158676
rect 343652 158612 343653 158676
rect 343587 158611 343653 158612
rect 343955 158676 344021 158677
rect 343955 158612 343956 158676
rect 344020 158612 344021 158676
rect 343955 158611 344021 158612
rect 342851 157996 342917 157997
rect 342851 157932 342852 157996
rect 342916 157932 342917 157996
rect 342851 157931 342917 157932
rect 341747 157860 341813 157861
rect 341747 157796 341748 157860
rect 341812 157796 341813 157860
rect 341747 157795 341813 157796
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 129454 344414 158000
rect 345246 157861 345306 159430
rect 345982 158677 346042 159430
rect 346350 159430 346444 159490
rect 347608 159490 347668 160106
rect 348288 159901 348348 160106
rect 348285 159900 348351 159901
rect 348285 159836 348286 159900
rect 348350 159836 348351 159900
rect 348285 159835 348351 159836
rect 348696 159490 348756 160106
rect 349784 159490 349844 160106
rect 351008 159765 351068 160106
rect 351005 159764 351071 159765
rect 351005 159700 351006 159764
rect 351070 159700 351071 159764
rect 351005 159699 351071 159700
rect 351144 159490 351204 160106
rect 347608 159430 347698 159490
rect 348696 159430 348802 159490
rect 349784 159430 349906 159490
rect 345979 158676 346045 158677
rect 345979 158612 345980 158676
rect 346044 158612 346045 158676
rect 345979 158611 346045 158612
rect 346350 157861 346410 159430
rect 347638 157997 347698 159430
rect 348742 158677 348802 159430
rect 348739 158676 348805 158677
rect 348739 158612 348740 158676
rect 348804 158612 348805 158676
rect 348739 158611 348805 158612
rect 347635 157996 347701 157997
rect 347635 157932 347636 157996
rect 347700 157932 347701 157996
rect 347635 157931 347701 157932
rect 345243 157860 345309 157861
rect 345243 157796 345244 157860
rect 345308 157796 345309 157860
rect 345243 157795 345309 157796
rect 346347 157860 346413 157861
rect 346347 157796 346348 157860
rect 346412 157796 346413 157860
rect 346347 157795 346413 157796
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 133954 348914 158000
rect 349846 157453 349906 159430
rect 351134 159430 351204 159490
rect 352232 159490 352292 160106
rect 353320 159490 353380 160106
rect 353592 159765 353652 160106
rect 353589 159764 353655 159765
rect 353589 159700 353590 159764
rect 353654 159700 353655 159764
rect 353589 159699 353655 159700
rect 354408 159490 354468 160106
rect 355768 159490 355828 160106
rect 356040 159765 356100 160106
rect 356037 159764 356103 159765
rect 356037 159700 356038 159764
rect 356102 159700 356103 159764
rect 356037 159699 356103 159700
rect 352232 159430 352298 159490
rect 353320 159430 353402 159490
rect 354408 159430 354506 159490
rect 351134 157453 351194 159430
rect 352238 157453 352298 159430
rect 353342 158269 353402 159430
rect 353339 158268 353405 158269
rect 353339 158204 353340 158268
rect 353404 158204 353405 158268
rect 353339 158203 353405 158204
rect 349843 157452 349909 157453
rect 349843 157388 349844 157452
rect 349908 157388 349909 157452
rect 349843 157387 349909 157388
rect 351131 157452 351197 157453
rect 351131 157388 351132 157452
rect 351196 157388 351197 157452
rect 351131 157387 351197 157388
rect 352235 157452 352301 157453
rect 352235 157388 352236 157452
rect 352300 157388 352301 157452
rect 352235 157387 352301 157388
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 138454 353414 158000
rect 354446 157453 354506 159430
rect 355734 159430 355828 159490
rect 356992 159490 357052 160106
rect 358080 159490 358140 160106
rect 358488 159490 358548 160106
rect 359168 159490 359228 160106
rect 360936 159765 360996 160106
rect 363520 159901 363580 160106
rect 363517 159900 363583 159901
rect 363517 159836 363518 159900
rect 363582 159836 363583 159900
rect 363517 159835 363583 159836
rect 360933 159764 360999 159765
rect 360933 159700 360934 159764
rect 360998 159700 360999 159764
rect 360933 159699 360999 159700
rect 365968 159490 366028 160106
rect 368280 159490 368340 160106
rect 371000 159901 371060 160106
rect 370997 159900 371063 159901
rect 370997 159836 370998 159900
rect 371062 159836 371063 159900
rect 370997 159835 371063 159836
rect 373448 159490 373508 160106
rect 356992 159430 357082 159490
rect 358080 159430 358186 159490
rect 358488 159430 358554 159490
rect 359168 159430 359290 159490
rect 355734 158677 355794 159430
rect 357022 158677 357082 159430
rect 355731 158676 355797 158677
rect 355731 158612 355732 158676
rect 355796 158612 355797 158676
rect 355731 158611 355797 158612
rect 357019 158676 357085 158677
rect 357019 158612 357020 158676
rect 357084 158612 357085 158676
rect 357019 158611 357085 158612
rect 358126 158541 358186 159430
rect 358494 158677 358554 159430
rect 358491 158676 358557 158677
rect 358491 158612 358492 158676
rect 358556 158612 358557 158676
rect 358491 158611 358557 158612
rect 358123 158540 358189 158541
rect 358123 158476 358124 158540
rect 358188 158476 358189 158540
rect 358123 158475 358189 158476
rect 354443 157452 354509 157453
rect 354443 157388 354444 157452
rect 354508 157388 354509 157452
rect 354443 157387 354509 157388
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 142954 357914 158000
rect 359230 157589 359290 159430
rect 365854 159430 366028 159490
rect 368246 159430 368340 159490
rect 373398 159430 373508 159490
rect 375896 159490 375956 160106
rect 378480 159490 378540 160106
rect 380928 159490 380988 160106
rect 383512 159490 383572 160106
rect 385960 159490 386020 160106
rect 388544 159490 388604 160106
rect 375896 159430 376034 159490
rect 378480 159430 378610 159490
rect 380928 159430 381002 159490
rect 383512 159430 383578 159490
rect 365854 158677 365914 159430
rect 368246 158677 368306 159430
rect 373398 158677 373458 159430
rect 375974 158677 376034 159430
rect 378550 158677 378610 159430
rect 380942 158677 381002 159430
rect 383518 158677 383578 159430
rect 385910 159430 386020 159490
rect 388486 159430 388604 159490
rect 390992 159490 391052 160106
rect 393440 159490 393500 160106
rect 395888 159490 395948 160106
rect 398472 159490 398532 160106
rect 390992 159430 391122 159490
rect 393440 159430 393514 159490
rect 385910 158677 385970 159430
rect 388486 158677 388546 159430
rect 391062 158677 391122 159430
rect 393454 158677 393514 159430
rect 395846 159430 395948 159490
rect 398422 159430 398532 159490
rect 400920 159490 400980 160106
rect 403368 159490 403428 160106
rect 405952 159490 406012 160106
rect 400920 159430 401058 159490
rect 403368 159430 403450 159490
rect 405952 159430 406026 159490
rect 395846 158677 395906 159430
rect 398422 158677 398482 159430
rect 400998 158677 401058 159430
rect 403390 158677 403450 159430
rect 405966 158677 406026 159430
rect 365851 158676 365917 158677
rect 365851 158612 365852 158676
rect 365916 158612 365917 158676
rect 365851 158611 365917 158612
rect 368243 158676 368309 158677
rect 368243 158612 368244 158676
rect 368308 158612 368309 158676
rect 368243 158611 368309 158612
rect 373395 158676 373461 158677
rect 373395 158612 373396 158676
rect 373460 158612 373461 158676
rect 373395 158611 373461 158612
rect 375971 158676 376037 158677
rect 375971 158612 375972 158676
rect 376036 158612 376037 158676
rect 375971 158611 376037 158612
rect 378547 158676 378613 158677
rect 378547 158612 378548 158676
rect 378612 158612 378613 158676
rect 378547 158611 378613 158612
rect 380939 158676 381005 158677
rect 380939 158612 380940 158676
rect 381004 158612 381005 158676
rect 380939 158611 381005 158612
rect 383515 158676 383581 158677
rect 383515 158612 383516 158676
rect 383580 158612 383581 158676
rect 383515 158611 383581 158612
rect 385907 158676 385973 158677
rect 385907 158612 385908 158676
rect 385972 158612 385973 158676
rect 385907 158611 385973 158612
rect 388483 158676 388549 158677
rect 388483 158612 388484 158676
rect 388548 158612 388549 158676
rect 388483 158611 388549 158612
rect 391059 158676 391125 158677
rect 391059 158612 391060 158676
rect 391124 158612 391125 158676
rect 391059 158611 391125 158612
rect 393451 158676 393517 158677
rect 393451 158612 393452 158676
rect 393516 158612 393517 158676
rect 393451 158611 393517 158612
rect 395843 158676 395909 158677
rect 395843 158612 395844 158676
rect 395908 158612 395909 158676
rect 395843 158611 395909 158612
rect 398419 158676 398485 158677
rect 398419 158612 398420 158676
rect 398484 158612 398485 158676
rect 398419 158611 398485 158612
rect 400995 158676 401061 158677
rect 400995 158612 400996 158676
rect 401060 158612 401061 158676
rect 400995 158611 401061 158612
rect 403387 158676 403453 158677
rect 403387 158612 403388 158676
rect 403452 158612 403453 158676
rect 403387 158611 403453 158612
rect 405963 158676 406029 158677
rect 405963 158612 405964 158676
rect 406028 158612 406029 158676
rect 405963 158611 406029 158612
rect 359227 157588 359293 157589
rect 359227 157524 359228 157588
rect 359292 157524 359293 157588
rect 359227 157523 359293 157524
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 147454 362414 158000
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 151954 366914 158000
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 156454 371414 158000
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 124954 375914 158000
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 129454 380414 158000
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 133954 384914 158000
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 138454 389414 158000
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 142954 393914 158000
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 147454 398414 158000
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 151954 402914 158000
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 156454 407414 158000
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 124954 411914 158000
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 129454 416414 158000
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 133954 420914 158000
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 138454 425414 158000
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 142954 429914 158000
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 147454 434414 158000
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 437430 3637 437490 297331
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 439083 261492 439149 261493
rect 439083 261428 439084 261492
rect 439148 261428 439149 261492
rect 439083 261427 439149 261428
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 437611 248300 437677 248301
rect 437611 248236 437612 248300
rect 437676 248236 437677 248300
rect 437611 248235 437677 248236
rect 437427 3636 437493 3637
rect 437427 3572 437428 3636
rect 437492 3572 437493 3636
rect 437427 3571 437493 3572
rect 437614 3501 437674 248235
rect 437795 245308 437861 245309
rect 438294 245308 438914 259398
rect 437795 245244 437796 245308
rect 437860 245244 437861 245308
rect 437795 245243 437861 245244
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 437611 3500 437677 3501
rect 437611 3436 437612 3500
rect 437676 3436 437677 3500
rect 437611 3435 437677 3436
rect 437798 3365 437858 245243
rect 438294 151954 438914 158000
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 437795 3364 437861 3365
rect 437795 3300 437796 3364
rect 437860 3300 437861 3364
rect 437795 3299 437861 3300
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 -1306 438914 7398
rect 439086 3501 439146 261427
rect 439454 71909 439514 444347
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 439451 71908 439517 71909
rect 439451 71844 439452 71908
rect 439516 71844 439517 71908
rect 439451 71843 439517 71844
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 439083 3500 439149 3501
rect 439083 3436 439084 3500
rect 439148 3436 439149 3500
rect 439083 3435 439149 3436
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< obsm4 >>
rect 220000 547986 356620 563308
rect 220000 547366 220272 547986
rect 220620 547366 356000 547986
rect 356348 547366 356620 547986
rect 220000 543486 356620 547366
rect 220000 542866 220952 543486
rect 221300 542866 355320 543486
rect 355668 542866 356620 543486
rect 220000 511986 356620 542866
rect 220000 511366 220272 511986
rect 220620 511366 356000 511986
rect 356348 511366 356620 511986
rect 220000 507486 356620 511366
rect 220000 506866 220952 507486
rect 221300 506866 355320 507486
rect 355668 506866 356620 507486
rect 220000 480080 356620 506866
rect 220000 480000 236056 480080
rect 236116 480000 237144 480080
rect 237204 480000 238232 480080
rect 238292 480000 239592 480080
rect 239652 480000 240544 480080
rect 240604 480000 241768 480080
rect 241828 480000 243128 480080
rect 243188 480000 244216 480080
rect 244276 480000 245440 480080
rect 245500 480000 246528 480080
rect 246588 480000 247616 480080
rect 247676 480000 248296 480080
rect 248356 480000 248704 480080
rect 248764 480000 250064 480080
rect 250124 480000 250744 480080
rect 250804 480000 251288 480080
rect 251348 480000 252376 480080
rect 252436 480000 253464 480080
rect 253524 480000 253600 480080
rect 253660 480000 254552 480080
rect 254612 480000 255912 480080
rect 255972 480000 256048 480080
rect 256108 480000 257000 480080
rect 257060 480000 258088 480080
rect 258148 480000 258496 480080
rect 258556 480000 259448 480080
rect 259508 480000 260672 480080
rect 260732 480000 261080 480080
rect 261140 480000 261760 480080
rect 261820 480000 262848 480080
rect 262908 480000 263528 480080
rect 263588 480000 263936 480080
rect 263996 480000 265296 480080
rect 265356 480000 265976 480080
rect 266036 480000 266384 480080
rect 266444 480000 267608 480080
rect 267668 480000 268288 480080
rect 268348 480000 268696 480080
rect 268756 480000 269784 480080
rect 269844 480000 271008 480080
rect 271068 480000 271144 480080
rect 271204 480000 272232 480080
rect 272292 480000 273320 480080
rect 273380 480000 273592 480080
rect 273652 480000 274408 480080
rect 274468 480000 275768 480080
rect 275828 480000 276040 480080
rect 276100 480000 276992 480080
rect 277052 480000 278080 480080
rect 278140 480000 278488 480080
rect 278548 480000 279168 480080
rect 279228 480000 280936 480080
rect 280996 480000 283520 480080
rect 283580 480000 285968 480080
rect 286028 480000 288280 480080
rect 288340 480000 291000 480080
rect 291060 480000 293448 480080
rect 293508 480000 295896 480080
rect 295956 480000 298480 480080
rect 298540 480000 300928 480080
rect 300988 480000 303512 480080
rect 303572 480000 305960 480080
rect 306020 480000 308544 480080
rect 308604 480000 310992 480080
rect 311052 480000 313440 480080
rect 313500 480000 315888 480080
rect 315948 480000 318472 480080
rect 318532 480000 320920 480080
rect 320980 480000 323368 480080
rect 323428 480000 325952 480080
rect 326012 480000 356620 480080
rect 100000 223986 236620 243308
rect 100000 223366 100272 223986
rect 100620 223366 236000 223986
rect 236348 223366 236620 223986
rect 100000 219486 236620 223366
rect 100000 218866 100952 219486
rect 101300 218866 235320 219486
rect 235668 218866 236620 219486
rect 100000 187986 236620 218866
rect 100000 187366 100272 187986
rect 100620 187366 236000 187986
rect 236348 187366 236620 187986
rect 100000 183486 236620 187366
rect 100000 182866 100952 183486
rect 101300 182866 235320 183486
rect 235668 182866 236620 183486
rect 100000 160106 236620 182866
rect 100000 160000 116056 160106
rect 116116 160000 117144 160106
rect 117204 160000 118232 160106
rect 118292 160000 119592 160106
rect 119652 160000 120544 160106
rect 120604 160000 121768 160106
rect 121828 160000 123128 160106
rect 123188 160000 124216 160106
rect 124276 160000 125440 160106
rect 125500 160000 126528 160106
rect 126588 160000 127616 160106
rect 127676 160000 128296 160106
rect 128356 160000 128704 160106
rect 128764 160000 130064 160106
rect 130124 160000 130744 160106
rect 130804 160000 131288 160106
rect 131348 160000 132376 160106
rect 132436 160000 133464 160106
rect 133524 160000 133600 160106
rect 133660 160000 134552 160106
rect 134612 160000 135912 160106
rect 135972 160000 136048 160106
rect 136108 160000 137000 160106
rect 137060 160000 138088 160106
rect 138148 160000 138496 160106
rect 138556 160000 139448 160106
rect 139508 160000 140672 160106
rect 140732 160000 141080 160106
rect 141140 160000 141760 160106
rect 141820 160000 142848 160106
rect 142908 160000 143528 160106
rect 143588 160000 143936 160106
rect 143996 160000 145296 160106
rect 145356 160000 145976 160106
rect 146036 160000 146384 160106
rect 146444 160000 147608 160106
rect 147668 160000 148288 160106
rect 148348 160000 148696 160106
rect 148756 160000 149784 160106
rect 149844 160000 151008 160106
rect 151068 160000 151144 160106
rect 151204 160000 152232 160106
rect 152292 160000 153320 160106
rect 153380 160000 153592 160106
rect 153652 160000 154408 160106
rect 154468 160000 155768 160106
rect 155828 160000 156040 160106
rect 156100 160000 156992 160106
rect 157052 160000 158080 160106
rect 158140 160000 158488 160106
rect 158548 160000 159168 160106
rect 159228 160000 160936 160106
rect 160996 160000 163520 160106
rect 163580 160000 165968 160106
rect 166028 160000 168280 160106
rect 168340 160000 171000 160106
rect 171060 160000 173448 160106
rect 173508 160000 175896 160106
rect 175956 160000 178480 160106
rect 178540 160000 180928 160106
rect 180988 160000 183512 160106
rect 183572 160000 185960 160106
rect 186020 160000 188544 160106
rect 188604 160000 190992 160106
rect 191052 160000 193440 160106
rect 193500 160000 195888 160106
rect 195948 160000 198472 160106
rect 198532 160000 200920 160106
rect 200980 160000 203368 160106
rect 203428 160000 205952 160106
rect 206012 160000 236620 160106
rect 300000 223986 436620 243308
rect 300000 223366 300272 223986
rect 300620 223366 436000 223986
rect 436348 223366 436620 223986
rect 300000 219486 436620 223366
rect 300000 218866 300952 219486
rect 301300 218866 435320 219486
rect 435668 218866 436620 219486
rect 300000 187986 436620 218866
rect 300000 187366 300272 187986
rect 300620 187366 436000 187986
rect 436348 187366 436620 187986
rect 300000 183486 436620 187366
rect 300000 182866 300952 183486
rect 301300 182866 435320 183486
rect 435668 182866 436620 183486
rect 300000 160106 436620 182866
rect 300000 160000 316056 160106
rect 316116 160000 317144 160106
rect 317204 160000 318232 160106
rect 318292 160000 319592 160106
rect 319652 160000 320544 160106
rect 320604 160000 321768 160106
rect 321828 160000 323128 160106
rect 323188 160000 324216 160106
rect 324276 160000 325440 160106
rect 325500 160000 326528 160106
rect 326588 160000 327616 160106
rect 327676 160000 328296 160106
rect 328356 160000 328704 160106
rect 328764 160000 330064 160106
rect 330124 160000 330744 160106
rect 330804 160000 331288 160106
rect 331348 160000 332376 160106
rect 332436 160000 333464 160106
rect 333524 160000 333600 160106
rect 333660 160000 334552 160106
rect 334612 160000 335912 160106
rect 335972 160000 336048 160106
rect 336108 160000 337000 160106
rect 337060 160000 338088 160106
rect 338148 160000 338496 160106
rect 338556 160000 339448 160106
rect 339508 160000 340672 160106
rect 340732 160000 341080 160106
rect 341140 160000 341760 160106
rect 341820 160000 342848 160106
rect 342908 160000 343528 160106
rect 343588 160000 343936 160106
rect 343996 160000 345296 160106
rect 345356 160000 345976 160106
rect 346036 160000 346384 160106
rect 346444 160000 347608 160106
rect 347668 160000 348288 160106
rect 348348 160000 348696 160106
rect 348756 160000 349784 160106
rect 349844 160000 351008 160106
rect 351068 160000 351144 160106
rect 351204 160000 352232 160106
rect 352292 160000 353320 160106
rect 353380 160000 353592 160106
rect 353652 160000 354408 160106
rect 354468 160000 355768 160106
rect 355828 160000 356040 160106
rect 356100 160000 356992 160106
rect 357052 160000 358080 160106
rect 358140 160000 358488 160106
rect 358548 160000 359168 160106
rect 359228 160000 360936 160106
rect 360996 160000 363520 160106
rect 363580 160000 365968 160106
rect 366028 160000 368280 160106
rect 368340 160000 371000 160106
rect 371060 160000 373448 160106
rect 373508 160000 375896 160106
rect 375956 160000 378480 160106
rect 378540 160000 380928 160106
rect 380988 160000 383512 160106
rect 383572 160000 385960 160106
rect 386020 160000 388544 160106
rect 388604 160000 390992 160106
rect 391052 160000 393440 160106
rect 393500 160000 395888 160106
rect 395948 160000 398472 160106
rect 398532 160000 400920 160106
rect 400980 160000 403368 160106
rect 403428 160000 405952 160106
rect 406012 160000 436620 160106
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 220328 547718 220564 547954
rect 220328 547398 220564 547634
rect 356056 547718 356292 547954
rect 356056 547398 356292 547634
rect 221008 543218 221244 543454
rect 221008 542898 221244 543134
rect 355376 543218 355612 543454
rect 355376 542898 355612 543134
rect 220328 511718 220564 511954
rect 220328 511398 220564 511634
rect 356056 511718 356292 511954
rect 356056 511398 356292 511634
rect 221008 507218 221244 507454
rect 221008 506898 221244 507134
rect 355376 507218 355612 507454
rect 355376 506898 355612 507134
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 249610 439718 249846 439954
rect 249610 439398 249846 439634
rect 280330 439718 280566 439954
rect 280330 439398 280566 439634
rect 311050 439718 311286 439954
rect 311050 439398 311286 439634
rect 341770 439718 342006 439954
rect 341770 439398 342006 439634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 234250 435218 234486 435454
rect 234250 434898 234486 435134
rect 264970 435218 265206 435454
rect 264970 434898 265206 435134
rect 295690 435218 295926 435454
rect 295690 434898 295926 435134
rect 326410 435218 326646 435454
rect 326410 434898 326646 435134
rect 357130 435218 357366 435454
rect 357130 434898 357366 435134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 249610 403718 249846 403954
rect 249610 403398 249846 403634
rect 280330 403718 280566 403954
rect 280330 403398 280566 403634
rect 311050 403718 311286 403954
rect 311050 403398 311286 403634
rect 341770 403718 342006 403954
rect 341770 403398 342006 403634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 234250 399218 234486 399454
rect 234250 398898 234486 399134
rect 264970 399218 265206 399454
rect 264970 398898 265206 399134
rect 295690 399218 295926 399454
rect 295690 398898 295926 399134
rect 326410 399218 326646 399454
rect 326410 398898 326646 399134
rect 357130 399218 357366 399454
rect 357130 398898 357366 399134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 249610 367718 249846 367954
rect 249610 367398 249846 367634
rect 280330 367718 280566 367954
rect 280330 367398 280566 367634
rect 311050 367718 311286 367954
rect 311050 367398 311286 367634
rect 341770 367718 342006 367954
rect 341770 367398 342006 367634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 234250 363218 234486 363454
rect 234250 362898 234486 363134
rect 264970 363218 265206 363454
rect 264970 362898 265206 363134
rect 295690 363218 295926 363454
rect 295690 362898 295926 363134
rect 326410 363218 326646 363454
rect 326410 362898 326646 363134
rect 357130 363218 357366 363454
rect 357130 362898 357366 363134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 249610 331718 249846 331954
rect 249610 331398 249846 331634
rect 280330 331718 280566 331954
rect 280330 331398 280566 331634
rect 311050 331718 311286 331954
rect 311050 331398 311286 331634
rect 341770 331718 342006 331954
rect 341770 331398 342006 331634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 234250 327218 234486 327454
rect 234250 326898 234486 327134
rect 264970 327218 265206 327454
rect 264970 326898 265206 327134
rect 295690 327218 295926 327454
rect 295690 326898 295926 327134
rect 326410 327218 326646 327454
rect 326410 326898 326646 327134
rect 357130 327218 357366 327454
rect 357130 326898 357366 327134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 100328 223718 100564 223954
rect 100328 223398 100564 223634
rect 236056 223718 236292 223954
rect 236056 223398 236292 223634
rect 101008 219218 101244 219454
rect 101008 218898 101244 219134
rect 235376 219218 235612 219454
rect 235376 218898 235612 219134
rect 100328 187718 100564 187954
rect 100328 187398 100564 187634
rect 236056 187718 236292 187954
rect 236056 187398 236292 187634
rect 101008 183218 101244 183454
rect 101008 182898 101244 183134
rect 235376 183218 235612 183454
rect 235376 182898 235612 183134
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 120218 119062 120454
rect 119146 120218 119382 120454
rect 118826 119898 119062 120134
rect 119146 119898 119382 120134
rect 118826 84218 119062 84454
rect 119146 84218 119382 84454
rect 118826 83898 119062 84134
rect 119146 83898 119382 84134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 124718 123562 124954
rect 123646 124718 123882 124954
rect 123326 124398 123562 124634
rect 123646 124398 123882 124634
rect 123326 88718 123562 88954
rect 123646 88718 123882 88954
rect 123326 88398 123562 88634
rect 123646 88398 123882 88634
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 133718 132562 133954
rect 132646 133718 132882 133954
rect 132326 133398 132562 133634
rect 132646 133398 132882 133634
rect 132326 97718 132562 97954
rect 132646 97718 132882 97954
rect 132326 97398 132562 97634
rect 132646 97398 132882 97634
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 138218 137062 138454
rect 137146 138218 137382 138454
rect 136826 137898 137062 138134
rect 137146 137898 137382 138134
rect 136826 102218 137062 102454
rect 137146 102218 137382 102454
rect 136826 101898 137062 102134
rect 137146 101898 137382 102134
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 106718 141562 106954
rect 141646 106718 141882 106954
rect 141326 106398 141562 106634
rect 141646 106398 141882 106634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 150326 115718 150562 115954
rect 150646 115718 150882 115954
rect 150326 115398 150562 115634
rect 150646 115398 150882 115634
rect 150326 79718 150562 79954
rect 150646 79718 150882 79954
rect 150326 79398 150562 79634
rect 150646 79398 150882 79634
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154826 120218 155062 120454
rect 155146 120218 155382 120454
rect 154826 119898 155062 120134
rect 155146 119898 155382 120134
rect 154826 84218 155062 84454
rect 155146 84218 155382 84454
rect 154826 83898 155062 84134
rect 155146 83898 155382 84134
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 124718 159562 124954
rect 159646 124718 159882 124954
rect 159326 124398 159562 124634
rect 159646 124398 159882 124634
rect 159326 88718 159562 88954
rect 159646 88718 159882 88954
rect 159326 88398 159562 88634
rect 159646 88398 159882 88634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 133718 168562 133954
rect 168646 133718 168882 133954
rect 168326 133398 168562 133634
rect 168646 133398 168882 133634
rect 168326 97718 168562 97954
rect 168646 97718 168882 97954
rect 168326 97398 168562 97634
rect 168646 97398 168882 97634
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 138218 173062 138454
rect 173146 138218 173382 138454
rect 172826 137898 173062 138134
rect 173146 137898 173382 138134
rect 172826 102218 173062 102454
rect 173146 102218 173382 102454
rect 172826 101898 173062 102134
rect 173146 101898 173382 102134
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 106718 177562 106954
rect 177646 106718 177882 106954
rect 177326 106398 177562 106634
rect 177646 106398 177882 106634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 186326 115718 186562 115954
rect 186646 115718 186882 115954
rect 186326 115398 186562 115634
rect 186646 115398 186882 115634
rect 186326 79718 186562 79954
rect 186646 79718 186882 79954
rect 186326 79398 186562 79634
rect 186646 79398 186882 79634
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 190826 120218 191062 120454
rect 191146 120218 191382 120454
rect 190826 119898 191062 120134
rect 191146 119898 191382 120134
rect 190826 84218 191062 84454
rect 191146 84218 191382 84454
rect 190826 83898 191062 84134
rect 191146 83898 191382 84134
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 300328 223718 300564 223954
rect 300328 223398 300564 223634
rect 436056 223718 436292 223954
rect 436056 223398 436292 223634
rect 301008 219218 301244 219454
rect 301008 218898 301244 219134
rect 435376 219218 435612 219454
rect 435376 218898 435612 219134
rect 300328 187718 300564 187954
rect 300328 187398 300564 187634
rect 436056 187718 436292 187954
rect 436056 187398 436292 187634
rect 301008 183218 301244 183454
rect 301008 182898 301244 183134
rect 435376 183218 435612 183454
rect 435376 182898 435612 183134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 220328 547954
rect 220564 547718 356056 547954
rect 356292 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 220328 547634
rect 220564 547398 356056 547634
rect 356292 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 221008 543454
rect 221244 543218 355376 543454
rect 355612 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 221008 543134
rect 221244 542898 355376 543134
rect 355612 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 220328 511954
rect 220564 511718 356056 511954
rect 356292 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 220328 511634
rect 220564 511398 356056 511634
rect 356292 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 221008 507454
rect 221244 507218 355376 507454
rect 355612 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 221008 507134
rect 221244 506898 355376 507134
rect 355612 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 249610 439954
rect 249846 439718 280330 439954
rect 280566 439718 311050 439954
rect 311286 439718 341770 439954
rect 342006 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 249610 439634
rect 249846 439398 280330 439634
rect 280566 439398 311050 439634
rect 311286 439398 341770 439634
rect 342006 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 234250 435454
rect 234486 435218 264970 435454
rect 265206 435218 295690 435454
rect 295926 435218 326410 435454
rect 326646 435218 357130 435454
rect 357366 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 234250 435134
rect 234486 434898 264970 435134
rect 265206 434898 295690 435134
rect 295926 434898 326410 435134
rect 326646 434898 357130 435134
rect 357366 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 249610 403954
rect 249846 403718 280330 403954
rect 280566 403718 311050 403954
rect 311286 403718 341770 403954
rect 342006 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 249610 403634
rect 249846 403398 280330 403634
rect 280566 403398 311050 403634
rect 311286 403398 341770 403634
rect 342006 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 234250 399454
rect 234486 399218 264970 399454
rect 265206 399218 295690 399454
rect 295926 399218 326410 399454
rect 326646 399218 357130 399454
rect 357366 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 234250 399134
rect 234486 398898 264970 399134
rect 265206 398898 295690 399134
rect 295926 398898 326410 399134
rect 326646 398898 357130 399134
rect 357366 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 249610 367954
rect 249846 367718 280330 367954
rect 280566 367718 311050 367954
rect 311286 367718 341770 367954
rect 342006 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 249610 367634
rect 249846 367398 280330 367634
rect 280566 367398 311050 367634
rect 311286 367398 341770 367634
rect 342006 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 234250 363454
rect 234486 363218 264970 363454
rect 265206 363218 295690 363454
rect 295926 363218 326410 363454
rect 326646 363218 357130 363454
rect 357366 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 234250 363134
rect 234486 362898 264970 363134
rect 265206 362898 295690 363134
rect 295926 362898 326410 363134
rect 326646 362898 357130 363134
rect 357366 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 249610 331954
rect 249846 331718 280330 331954
rect 280566 331718 311050 331954
rect 311286 331718 341770 331954
rect 342006 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 249610 331634
rect 249846 331398 280330 331634
rect 280566 331398 311050 331634
rect 311286 331398 341770 331634
rect 342006 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 234250 327454
rect 234486 327218 264970 327454
rect 265206 327218 295690 327454
rect 295926 327218 326410 327454
rect 326646 327218 357130 327454
rect 357366 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 234250 327134
rect 234486 326898 264970 327134
rect 265206 326898 295690 327134
rect 295926 326898 326410 327134
rect 326646 326898 357130 327134
rect 357366 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 100328 223954
rect 100564 223718 236056 223954
rect 236292 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 300328 223954
rect 300564 223718 436056 223954
rect 436292 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 100328 223634
rect 100564 223398 236056 223634
rect 236292 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 300328 223634
rect 300564 223398 436056 223634
rect 436292 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 101008 219454
rect 101244 219218 235376 219454
rect 235612 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 301008 219454
rect 301244 219218 435376 219454
rect 435612 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 101008 219134
rect 101244 218898 235376 219134
rect 235612 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 301008 219134
rect 301244 218898 435376 219134
rect 435612 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 100328 187954
rect 100564 187718 236056 187954
rect 236292 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 300328 187954
rect 300564 187718 436056 187954
rect 436292 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 100328 187634
rect 100564 187398 236056 187634
rect 236292 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 300328 187634
rect 300564 187398 436056 187634
rect 436292 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 101008 183454
rect 101244 183218 235376 183454
rect 235612 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 301008 183454
rect 301244 183218 435376 183454
rect 435612 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 101008 183134
rect 101244 182898 235376 183134
rect 235612 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 301008 183134
rect 301244 182898 435376 183134
rect 435612 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 136826 138454
rect 137062 138218 137146 138454
rect 137382 138218 172826 138454
rect 173062 138218 173146 138454
rect 173382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 136826 138134
rect 137062 137898 137146 138134
rect 137382 137898 172826 138134
rect 173062 137898 173146 138134
rect 173382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 132326 133954
rect 132562 133718 132646 133954
rect 132882 133718 168326 133954
rect 168562 133718 168646 133954
rect 168882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 132326 133634
rect 132562 133398 132646 133634
rect 132882 133398 168326 133634
rect 168562 133398 168646 133634
rect 168882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 123326 124954
rect 123562 124718 123646 124954
rect 123882 124718 159326 124954
rect 159562 124718 159646 124954
rect 159882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 123326 124634
rect 123562 124398 123646 124634
rect 123882 124398 159326 124634
rect 159562 124398 159646 124634
rect 159882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 118826 120454
rect 119062 120218 119146 120454
rect 119382 120218 154826 120454
rect 155062 120218 155146 120454
rect 155382 120218 190826 120454
rect 191062 120218 191146 120454
rect 191382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 118826 120134
rect 119062 119898 119146 120134
rect 119382 119898 154826 120134
rect 155062 119898 155146 120134
rect 155382 119898 190826 120134
rect 191062 119898 191146 120134
rect 191382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 150326 115954
rect 150562 115718 150646 115954
rect 150882 115718 186326 115954
rect 186562 115718 186646 115954
rect 186882 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 150326 115634
rect 150562 115398 150646 115634
rect 150882 115398 186326 115634
rect 186562 115398 186646 115634
rect 186882 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 141326 106954
rect 141562 106718 141646 106954
rect 141882 106718 177326 106954
rect 177562 106718 177646 106954
rect 177882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 141326 106634
rect 141562 106398 141646 106634
rect 141882 106398 177326 106634
rect 177562 106398 177646 106634
rect 177882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 136826 102454
rect 137062 102218 137146 102454
rect 137382 102218 172826 102454
rect 173062 102218 173146 102454
rect 173382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 136826 102134
rect 137062 101898 137146 102134
rect 137382 101898 172826 102134
rect 173062 101898 173146 102134
rect 173382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 132326 97954
rect 132562 97718 132646 97954
rect 132882 97718 168326 97954
rect 168562 97718 168646 97954
rect 168882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 132326 97634
rect 132562 97398 132646 97634
rect 132882 97398 168326 97634
rect 168562 97398 168646 97634
rect 168882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 123326 88954
rect 123562 88718 123646 88954
rect 123882 88718 159326 88954
rect 159562 88718 159646 88954
rect 159882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 123326 88634
rect 123562 88398 123646 88634
rect 123882 88398 159326 88634
rect 159562 88398 159646 88634
rect 159882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 118826 84454
rect 119062 84218 119146 84454
rect 119382 84218 154826 84454
rect 155062 84218 155146 84454
rect 155382 84218 190826 84454
rect 191062 84218 191146 84454
rect 191382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 118826 84134
rect 119062 83898 119146 84134
rect 119382 83898 154826 84134
rect 155062 83898 155146 84134
rect 155382 83898 190826 84134
rect 191062 83898 191146 84134
rect 191382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 150326 79954
rect 150562 79718 150646 79954
rect 150882 79718 186326 79954
rect 186562 79718 186646 79954
rect 186882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 150326 79634
rect 150562 79398 150646 79634
rect 150882 79398 186326 79634
rect 186562 79398 186646 79634
rect 186882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
<< obsm5 >>
rect 0 700986 584000 704000
rect 0 696486 584000 700366
rect 0 691986 584000 695866
rect 0 687486 584000 691366
rect 0 682986 584000 686866
rect 0 678486 584000 682366
rect 0 673986 584000 677866
rect 0 669486 584000 673366
rect 0 664986 584000 668866
rect 0 660486 584000 664366
rect 0 655986 584000 659866
rect 0 651486 584000 655366
rect 0 646986 584000 650866
rect 0 642486 584000 646366
rect 0 637986 584000 641866
rect 0 633486 584000 637366
rect 0 628986 584000 632866
rect 0 624486 584000 628366
rect 0 619986 584000 623866
rect 0 615486 584000 619366
rect 0 610986 584000 614866
rect 0 606486 584000 610366
rect 0 601986 584000 605866
rect 0 597486 584000 601366
rect 0 592986 584000 596866
rect 0 588486 584000 592366
rect 0 583986 584000 587866
rect 0 579486 584000 583366
rect 0 574986 584000 578866
rect 0 570486 584000 574366
rect 0 565986 584000 569866
rect 0 561486 584000 565366
rect 0 556986 584000 560866
rect 0 552486 584000 556366
rect 0 547986 584000 551866
rect 0 543486 584000 547366
rect 0 538986 584000 542866
rect 0 534486 584000 538366
rect 0 529986 584000 533866
rect 0 525486 584000 529366
rect 0 520986 584000 524866
rect 0 516486 584000 520366
rect 0 511986 584000 515866
rect 0 507486 584000 511366
rect 0 502986 584000 506866
rect 0 498486 584000 502366
rect 0 493986 584000 497866
rect 0 489486 584000 493366
rect 0 484986 584000 488866
rect 0 480486 584000 484366
rect 0 475986 584000 479866
rect 0 471486 584000 475366
rect 0 466986 584000 470866
rect 0 462486 584000 466366
rect 0 457986 584000 461866
rect 0 453486 584000 457366
rect 0 448986 584000 452866
rect 0 444486 584000 448366
rect 0 439986 584000 443866
rect 0 435486 584000 439366
rect 0 430986 584000 434866
rect 0 426486 584000 430366
rect 0 421986 584000 425866
rect 0 417486 584000 421366
rect 0 412986 584000 416866
rect 0 408486 584000 412366
rect 0 403986 584000 407866
rect 0 399486 584000 403366
rect 0 394986 584000 398866
rect 0 390486 584000 394366
rect 0 385986 584000 389866
rect 0 381486 584000 385366
rect 0 376986 584000 380866
rect 0 372486 584000 376366
rect 0 367986 584000 371866
rect 0 363486 584000 367366
rect 0 358986 584000 362866
rect 0 354486 584000 358366
rect 0 349986 584000 353866
rect 0 345486 584000 349366
rect 0 340986 584000 344866
rect 0 336486 584000 340366
rect 0 331986 584000 335866
rect 0 327486 584000 331366
rect 0 322986 584000 326866
rect 0 318486 584000 322366
rect 0 313986 584000 317866
rect 0 309486 584000 313366
rect 0 304986 584000 308866
rect 0 300486 584000 304366
rect 0 295986 584000 299866
rect 0 291486 584000 295366
rect 0 286986 584000 290866
rect 0 282486 584000 286366
rect 0 277986 584000 281866
rect 0 273486 584000 277366
rect 0 268986 584000 272866
rect 0 264486 584000 268366
rect 0 259986 584000 263866
rect 0 255486 584000 259366
rect 0 250986 584000 254866
rect 0 246486 584000 250366
rect 0 241986 584000 245866
rect 0 237486 584000 241366
rect 0 232986 584000 236866
rect 0 228486 584000 232366
rect 0 223986 584000 227866
rect 0 219486 584000 223366
rect 0 214986 584000 218866
rect 0 210486 584000 214366
rect 0 205986 584000 209866
rect 0 201486 584000 205366
rect 0 196986 584000 200866
rect 0 192486 584000 196366
rect 0 187986 584000 191866
rect 0 183486 584000 187366
rect 0 178986 584000 182866
rect 0 174486 584000 178366
rect 0 169986 584000 173866
rect 0 165486 584000 169366
rect 0 160986 584000 164866
rect 0 156486 584000 160366
rect 0 151986 584000 155866
rect 0 147486 584000 151366
rect 0 142986 584000 146866
rect 0 138486 584000 142366
rect 0 133986 584000 137866
rect 0 129486 584000 133366
rect 0 124986 584000 128866
rect 0 120486 584000 124366
rect 0 115986 584000 119866
rect 0 111486 584000 115366
rect 0 106986 584000 110866
rect 0 102486 584000 106366
rect 0 97986 584000 101866
rect 0 93486 584000 97366
rect 0 88986 584000 92866
rect 0 84486 584000 88366
rect 0 79986 584000 83866
rect 0 75486 584000 79366
rect 0 70986 584000 74866
rect 0 66486 584000 70366
rect 0 61986 584000 65866
rect 0 57486 584000 61366
rect 0 52986 584000 56866
rect 0 48486 584000 52366
rect 0 43986 584000 47866
rect 0 39486 584000 43366
rect 0 34986 584000 38866
rect 0 30486 584000 34366
rect 0 25986 584000 29866
rect 0 21486 584000 25366
rect 0 16986 584000 20866
rect 0 12486 584000 16366
rect 0 7986 584000 11866
rect 0 3486 584000 7366
rect 0 0 584000 2866
use sky130_sram_2kbyte_1rw1r_32x512_8  dram_inst
timestamp 0
transform 1 0 220000 0 1 480000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  iram_inst_A
timestamp 0
transform 1 0 100000 0 1 160000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  iram_inst_B
timestamp 0
transform 1 0 300000 0 1 160000
box 0 0 136620 83308
use rvj1_caravel_soc  rvj1_soc
timestamp 0
transform 1 0 230000 0 1 310400
box 1066 0 129758 133023
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 158000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 245308 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 158000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 245308 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 158000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 245308 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 158000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 245308 218414 478000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 565308 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 308400 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 565308 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 308400 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 565308 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 158000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 245308 326414 308400 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 565308 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 158000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 245308 362414 308400 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 445423 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 158000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 245308 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 158000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 245308 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 158000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 245308 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 158000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 245308 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 158000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 245308 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 158000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 245308 227414 478000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 565308 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 308400 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 565308 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 158000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 245308 299414 308400 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 565308 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 158000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 245308 335414 308400 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 565308 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 158000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 245308 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 158000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 245308 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 158000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 245308 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 158000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 245308 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 158000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 245308 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 158000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 565308 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 308400 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 565308 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 158000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 565308 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 158000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 565308 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 158000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 245308 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 158000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 245308 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 158000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 245308 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 158000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 245308 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 158000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 245308 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 158000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 245308 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 308400 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 565308 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 308400 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 565308 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 158000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 245308 317414 308400 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 565308 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 158000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 245308 353414 308400 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 565308 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 158000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 245308 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 158000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 245308 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 158000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 245308 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 158000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 245308 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 158000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 245308 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 308400 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 565308 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 308400 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 565308 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 158000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 565308 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 158000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 565308 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 158000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 245308 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 158000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 245308 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 158000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 245308 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 158000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 245308 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 158000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 245308 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 158000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 245308 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 308400 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 565308 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 308400 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 565308 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 158000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 245308 321914 308400 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 565308 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 158000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 245308 357914 308400 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 565308 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 158000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 245308 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 158000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 245308 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 158000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 245308 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 158000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 245308 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 158000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 245308 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 158000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 245308 222914 478000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 565308 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 308400 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 565308 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 308400 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 565308 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 158000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 245308 330914 308400 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 565308 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 158000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 245308 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 158000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 245308 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 158000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 245308 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 158000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 245308 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 158000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 245308 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 158000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 245308 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 158000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 245308 231914 308400 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 565308 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 308400 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 565308 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 158000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 245308 303914 308400 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 565308 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 158000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 245308 339914 308400 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 565308 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 158000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 245308 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 158000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 245308 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
